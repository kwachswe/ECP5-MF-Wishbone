
--
--------------------------------------------------------------------------------
--
-- File ID     : $Id: pcie_vhdl_test_case-pb.vhd 118 2022-01-17 23:26:12Z  $
-- Generated   : $LastChangedDate: 2022-01-18 00:26:12 +0100 (Tue, 18 Jan 2022) $
-- Revision    : $LastChangedRevision: 118 $
--
--------------------------------------------------------------------------------

Package Body pcie_vhdl_test_case_pkg is
   procedure run_test(signal clk : in    std_logic;
                      signal sv  : inout t_bfm_stim;
                      signal rv  : in    t_bfm_resp;
                             id  : in    natural := 0) is
   begin
      wait;
   end procedure; 

End pcie_vhdl_test_case_pkg;
