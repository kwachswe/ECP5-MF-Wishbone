module pcie_mfx1_top (
input wire ix_clk_125 ,
input wire [8 - 1 : 0] ix_dec_wb_cyc ,
input wire ix_ipx_dl_up ,
input wire ix_ipx_malf_tlp ,
input wire [16 - 1 : 0] ix_ipx_rx_data ,
input wire ix_ipx_rx_end ,
input wire ix_ipx_rx_st ,
input wire [12 : 0] ix_ipx_tx_ca_cpld ,
input wire [8 : 0] ix_ipx_tx_ca_cplh ,
input wire [12 : 0] ix_ipx_tx_ca_npd ,
input wire [8 : 0] ix_ipx_tx_ca_nph ,
input wire [12 : 0] ix_ipx_tx_ca_pd ,
input wire [8 : 0] ix_ipx_tx_ca_ph ,
input wire ix_ipx_tx_rdy ,
input wire [ 1 + 1 + 1 + 1 + 1 + 1 + 1 + 1 - 1 : 0] ix_pci_int_req ,
input wire ix_rst_n ,
input wire ix_wbm_ack ,
input wire [32 - 1 : 0] ix_wbm_dat ,
input wire [48 - 1 : 0] ix_wbs_adr ,
input wire [1 : 0] ix_wbs_bte ,
input wire [2 : 0] ix_wbs_cti ,
input wire [7 : 0] ix_wbs_cyc ,
input wire [32 - 1 : 0] ix_wbs_dat ,
input wire [(32 / 8) - 1 : 0] ix_wbs_sel ,
input wire ix_wbs_stb ,
input wire ix_wbs_we ,
output wire [16 - 1 : 0] ox_dec_adr ,
output wire [5 : 0] ox_dec_bar_hit ,
output wire [7 : 0] ox_dec_func_hit ,
output wire [7 : 0] ox_ipx_cc_npd_num ,
output wire [7 : 0] ox_ipx_cc_pd_num ,
output wire ox_ipx_cc_processed_npd ,
output wire ox_ipx_cc_processed_nph ,
output wire ox_ipx_cc_processed_pd ,
output wire ox_ipx_cc_processed_ph ,
output wire [16 - 1 : 0] ox_ipx_tx_data ,
output wire ox_ipx_tx_end ,
output wire ox_ipx_tx_req ,
output wire ox_ipx_tx_st ,
output wire [7 : 0] ox_sys_rst_func_n ,
output wire ox_sys_rst_n ,
output wire [16 - 1 : 0] ox_wbm_adr ,
output wire [1 : 0] ox_wbm_bte ,
output wire [2 : 0] ox_wbm_cti ,
output wire [8 - 1 : 0] ox_wbm_cyc ,
output wire [32 - 1 : 0] ox_wbm_dat ,
output wire [(32 / 8) - 1 : 0] ox_wbm_sel ,
output wire ox_wbm_stb ,
output wire ox_wbm_we ,
output wire ox_wbs_ack ,
output wire [32 - 1 : 0] ox_wbs_dat ,
output wire ox_wbs_err
   );
endmodule
