
//    
//    Copyright Ing. Buero Gardiner, 2007 - 2012
//     
//------------------------------------------------------------------------------
//
// File ID     : $Id: pcie_mfdev_v6.v 3810 2017-12-04 10:56:13Z  $
// Generated   : $LastChangedDate: 2017-12-04 11:56:13 +0100 (Mon, 04 Dec 2017) $
// Revision    : $LastChangedRevision: 3810 $
//
//------------------------------------------------------------------------------

`include "pci_exp_params.v" 
 
`timescale 1 ns / 1 ps
module credit_config (
   output wire          ox_fc_cpld_infinite,
   output wire          ox_fc_cplh_infinite,
   output wire          ox_fc_npd_infinite, 
   output wire          ox_fc_nph_infinite,
   output wire          ox_fc_pd_infinite,    
   output wire          ox_fc_ph_infinite,
   output wire [6:0]    ox_io_space_sel,
   output wire [7:0]    ox_hw_rev,
   output wire [15:0]   ox_subsys_id
   );

   wire [31:0]    w_init_reg_8;
   wire [31:0]    w_init_reg_2c;
      
   assign ox_fc_ph_infinite   = ( `INIT_PH_FC_VC0 == 0)   ? 1'b1 : 1'b0;
   assign ox_fc_pd_infinite   = ( `INIT_PD_FC_VC0 == 0)   ? 1'b1 : 1'b0;
   assign ox_fc_nph_infinite  = ( `INIT_NPH_FC_VC0 == 0)  ? 1'b1 : 1'b0;
   assign ox_fc_npd_infinite  = ( `INIT_NPD_FC_VC0 == 0)  ? 1'b1 : 1'b0;
   
   assign ox_io_space_sel[0]  = `INIT_REG_010 & 1'b1;
   assign ox_io_space_sel[1]  = `INIT_REG_014 & 1'b1;
   assign ox_io_space_sel[2]  = `INIT_REG_018 & 1'b1;
   assign ox_io_space_sel[3]  = `INIT_REG_01C & 1'b1;
   assign ox_io_space_sel[4]  = `INIT_REG_020 & 1'b1;
   assign ox_io_space_sel[5]  = `INIT_REG_024 & 1'b1;
   assign ox_io_space_sel[6]  = 1'b0;
   
   assign ox_hw_rev           = w_init_reg_8[7:0];
   
   assign ox_subsys_id        = w_init_reg_2c[31:16];
   
   `ifdef INIT_CPLH_FC_VC0
      assign ox_fc_cplh_infinite = ( `INIT_CPLH_FC_VC0 == 0) ? 1'b1 : 1'b0;
   `else
      assign ox_fc_cplh_infinite = 1'b1;
   `endif
   
   `ifdef INIT_CPLD_FC_VC0
      assign ox_fc_cpld_infinite = ( `INIT_CPLD_FC_VC0 == 0) ? 1'b1 : 1'b0;
   `else
      assign ox_fc_cpld_infinite = 1'b1;
   `endif
   
   assign w_init_reg_8  = `INIT_REG_008;
   assign w_init_reg_2c = `INIT_REG_02C;
   
endmodule
  `timescale 1 ns / 1 ps
module I6B46C5BDF6C2841AE2EEF22D18B3C8B9 # (parameter ID93CAA7BF31348EA47B29E962BD456C7 = 4, parameter IDD54D6BED81F43FAE3E38E047FDC453C
= 4, parameter I61D0345D311EC6FFC08DDDECE5F6127A = 256, parameter I5C6C6CD7723900C21B3A76E887CEE164 = 32, parameter
I64BB723AC8F87F7AEBA73BF190ED5F8F = 32, parameter I846B877ED5AEDADF389E2082E674F6A2 = 0 ) ( input wire ICCFB0F435B37370076102F325BC08D20 ,
input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire [I5C6C6CD7723900C21B3A76E887CEE164 + I846B877ED5AEDADF389E2082E674F6A2
- 1:0] I1A61D2CA45ECC28270C28826CD87FEC3 , input wire IC79EC9A9F373F4B71374BDF6EDD31DE6 , input wire I3DAC0A14B4001DD3A76D99313964C3AA ,
input wire IFF897FEF3F69926A750D8217ADD6AE1C , input wire I22B24791BA0E7AA2C686B1B2D776C636 , output wire [$clog2(I61D0345D311EC6FFC08DDDECE5F6127A )
- 1:0] I79D313D86841E5141E7629EA606D7AE9 , output wire I11CEFC90537A67CD1FF01400245362F2 , output wire [$clog2((I61D0345D311EC6FFC08DDDECE5F6127A
* (I5C6C6CD7723900C21B3A76E887CEE164 /I64BB723AC8F87F7AEBA73BF190ED5F8F )) + 1) - 1:0] ID7FCE45A65ADDB17F91F73A1B506BB5B ,
output wire [I64BB723AC8F87F7AEBA73BF190ED5F8F + I846B877ED5AEDADF389E2082E674F6A2 - 1:0] I125028C7446331521D0434C10E8B0007 ,
output wire I8BB939FF2AFDE7B2A1E480DCB61CE354 , output wire I41C63F948E534C7ED9F2471A44C922B2 , output wire I07E2A2E89C25B45C36871FC0931EC8EF ,
output wire [$clog2(I61D0345D311EC6FFC08DDDECE5F6127A ) - 1:0] I38B1AC532E13E69B05492C67EC7070BB , output wire I705C64753A50CDA034B5ACB332D71768 ,
output wire I102322A55721851004CB8E1F6AB50BDE , output wire [$clog2(I61D0345D311EC6FFC08DDDECE5F6127A + 1) - 1:0]
I233E0C0C8E5150F0CD8258F276D93942 , output wire IBE0D6810EBD63B5C428623C578CF6D3A , output wire I115E90220158F08B0465E99D7F2561D3
);  localparam ID4C318F5AC8B6BE2D0E1091653FE0983 = I5C6C6CD7723900C21B3A76E887CEE164 / I64BB723AC8F87F7AEBA73BF190ED5F8F ;
localparam I1AF585FFD3730CB75D8EA561C736B279 = ID93CAA7BF31348EA47B29E962BD456C7 ; localparam IB011AB9176BFCCD54AFA433401B9CC28
= ID93CAA7BF31348EA47B29E962BD456C7 + 1; localparam IC123CC1DD854BDF232C22DA342143DED = IDD54D6BED81F43FAE3E38E047FDC453C ;
localparam I41D54753579217A07881641483914F62 = IDD54D6BED81F43FAE3E38E047FDC453C + 1; localparam IEC3803494FB0D58F44099BF28643CCC0
= I5C6C6CD7723900C21B3A76E887CEE164 + I846B877ED5AEDADF389E2082E674F6A2 ; localparam IB7D40CABAAA60621C763075C02B43B42
= (ID4C318F5AC8B6BE2D0E1091653FE0983 == 1) ? ($clog2(ID4C318F5AC8B6BE2D0E1091653FE0983 ) + 1) : $clog2(ID4C318F5AC8B6BE2D0E1091653FE0983 );
localparam I2F6C1268D45752E3C34811C163B12775 = $clog2((I61D0345D311EC6FFC08DDDECE5F6127A * ID4C318F5AC8B6BE2D0E1091653FE0983 )
+ 1); localparam IAAE27A6B00F4178F2FC624379E618E64 = $clog2(I61D0345D311EC6FFC08DDDECE5F6127A + 1); localparam I2FB16649E1A7D4F99AB44B2AB26A8526
= $clog2(I61D0345D311EC6FFC08DDDECE5F6127A ); localparam ID5029CC947B009F8019DD7415E143367 = $clog2(I61D0345D311EC6FFC08DDDECE5F6127A
+ 1);  reg [IB7D40CABAAA60621C763075C02B43B42 - 1:0] I10F60E589450CD09FF7A498641DE26F8 ; reg [I2FB16649E1A7D4F99AB44B2AB26A8526
- 1:0] I3283453B42BD77672B8ACE724ACDA314 ; reg [I2FB16649E1A7D4F99AB44B2AB26A8526 - 1:0] IF8FA22381AE98928C01C1A8EF2CB0DC6 ;
reg I07E46217B3640C9CD06BF9B9D5D78F68 ; reg I7A2B537BEB4654059703B476744C6D18 ; reg I169F661B2921E0FA4AFB7C3794399862 ;
reg I87FD0B6E6C89D593796D3B1F631D5100 ; reg I4FD65DDA0EDE2F39B09EF91789B31572 ; reg [I2F6C1268D45752E3C34811C163B12775
- 1:0] IDDFF27981262750D43304A01A2EBF659 ; reg [I5C6C6CD7723900C21B3A76E887CEE164 + I846B877ED5AEDADF389E2082E674F6A2
- 1:0] I134B7C80786213E899F61495BA54C91C ; reg I00CE0BA4F77A2426865D797055E4C98A ; reg ID312B626B7C881C1A5210FC08BB95856 ;
reg I2E321486CBD81F71439B76F5D5BDCD93 ; reg [ID5029CC947B009F8019DD7415E143367 - 1:0] IDDCC249EE71726DC9EB38B3A433C91DB ;
reg I08DEC2092892554154AF13365E22F12A ; reg I6BE22F51BE43138B31F588DD2D062E1F ; reg I01F907CE74154BFFA0C1437099B21186 ;
reg [IAAE27A6B00F4178F2FC624379E618E64 - 1:0] IE1A203A1BCBBA5F947F638C3DFB65BF8 ; reg ID079750A1760FEED5898B26A23289BAD ;
reg I28ACD74043EE392893ABFA4360DDCD11 ; wire I38F39AED09C0507E780D3D35EA7FA06B ; wire I6316F5248B07D9065FBC7D67EDADC4EE ;
wire I2FAC1854542B2B806297DF5B4733F9D2 ; wire I61018042B0489325A4CD993FF565603E ;  assign I79D313D86841E5141E7629EA606D7AE9
= I3283453B42BD77672B8ACE724ACDA314 ; assign I11CEFC90537A67CD1FF01400245362F2 = I4FD65DDA0EDE2F39B09EF91789B31572 ;
assign ID7FCE45A65ADDB17F91F73A1B506BB5B = IDDFF27981262750D43304A01A2EBF659 ; assign I125028C7446331521D0434C10E8B0007
= (I846B877ED5AEDADF389E2082E674F6A2 == 0) ? I134B7C80786213E899F61495BA54C91C [I64BB723AC8F87F7AEBA73BF190ED5F8F
- 1:0] : {I134B7C80786213E899F61495BA54C91C [IEC3803494FB0D58F44099BF28643CCC0 - 1:I5C6C6CD7723900C21B3A76E887CEE164 ],
I134B7C80786213E899F61495BA54C91C [I64BB723AC8F87F7AEBA73BF190ED5F8F - 1:0]}; assign I8BB939FF2AFDE7B2A1E480DCB61CE354
= I00CE0BA4F77A2426865D797055E4C98A ; assign I41C63F948E534C7ED9F2471A44C922B2 = ID312B626B7C881C1A5210FC08BB95856 ;
assign I07E2A2E89C25B45C36871FC0931EC8EF = I2E321486CBD81F71439B76F5D5BDCD93 ; assign I38B1AC532E13E69B05492C67EC7070BB
= IF8FA22381AE98928C01C1A8EF2CB0DC6 ; assign I705C64753A50CDA034B5ACB332D71768 = I01F907CE74154BFFA0C1437099B21186 ;
assign I102322A55721851004CB8E1F6AB50BDE = I2FAC1854542B2B806297DF5B4733F9D2 ; assign I233E0C0C8E5150F0CD8258F276D93942
= IE1A203A1BCBBA5F947F638C3DFB65BF8 ; assign IBE0D6810EBD63B5C428623C578CF6D3A = ID079750A1760FEED5898B26A23289BAD ;
assign I115E90220158F08B0465E99D7F2561D3 = I28ACD74043EE392893ABFA4360DDCD11 ;  assign I38F39AED09C0507E780D3D35EA7FA06B
= (|I10F60E589450CD09FF7A498641DE26F8 ) ? 1'b0 : I6316F5248B07D9065FBC7D67EDADC4EE ; assign I6316F5248B07D9065FBC7D67EDADC4EE
= (I08DEC2092892554154AF13365E22F12A ) ? 1'b0 : (~I00CE0BA4F77A2426865D797055E4C98A | (|I10F60E589450CD09FF7A498641DE26F8 ));
assign I2FAC1854542B2B806297DF5B4733F9D2 = I22B24791BA0E7AA2C686B1B2D776C636 & ~ID079750A1760FEED5898B26A23289BAD ;
assign I61018042B0489325A4CD993FF565603E = (I6BE22F51BE43138B31F588DD2D062E1F ) ? 1'b0 : IFF897FEF3F69926A750D8217ADD6AE1C ;
 generate if (1'b1) begin : I50905559064282CED274D62360FCE175 reg [1:0] I102EDFAABB65014FC78C55AF4345F765 ; reg
[1:0] I69053399285CDFC39ECE32CB2CD079E5 ; reg [1:0] ICA80E74165E79AFA565A1A052BE49F09 ; task I8BE101CBEF6D2810BAC0C6F6AC8DA3B8 ;
begin I10F60E589450CD09FF7A498641DE26F8 <= {IB7D40CABAAA60621C763075C02B43B42 {1'b0}}; I3283453B42BD77672B8ACE724ACDA314
<= {I2FB16649E1A7D4F99AB44B2AB26A8526 {1'b0}}; IF8FA22381AE98928C01C1A8EF2CB0DC6 <= {I2FB16649E1A7D4F99AB44B2AB26A8526 {1'b0}};
I07E46217B3640C9CD06BF9B9D5D78F68 <= 1'b0; I7A2B537BEB4654059703B476744C6D18 <= 1'b0; I169F661B2921E0FA4AFB7C3794399862
<= 1'b0; I87FD0B6E6C89D593796D3B1F631D5100 <= 1'b0; I4FD65DDA0EDE2F39B09EF91789B31572 <= 1'b0; IDDFF27981262750D43304A01A2EBF659
<= {I2F6C1268D45752E3C34811C163B12775 {1'b0}}; I134B7C80786213E899F61495BA54C91C <= {IEC3803494FB0D58F44099BF28643CCC0 {1'b0}};
I00CE0BA4F77A2426865D797055E4C98A <= 1'b1; ID312B626B7C881C1A5210FC08BB95856 <= 1'b0; I2E321486CBD81F71439B76F5D5BDCD93
<= 1'b0; IDDCC249EE71726DC9EB38B3A433C91DB <= {ID5029CC947B009F8019DD7415E143367 {1'b0}}; I08DEC2092892554154AF13365E22F12A
<= 1'b1; I6BE22F51BE43138B31F588DD2D062E1F <= 1'b0; I01F907CE74154BFFA0C1437099B21186 <= 1'b0; IE1A203A1BCBBA5F947F638C3DFB65BF8
<= I61D0345D311EC6FFC08DDDECE5F6127A ; ID079750A1760FEED5898B26A23289BAD <= 1'b0; I28ACD74043EE392893ABFA4360DDCD11
<= 1'b0; end endtask always @(posedge ICCFB0F435B37370076102F325BC08D20 or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 )
begin if (I9ED2A9117D3AEAF54CBA7AD69083BCB7 == 1'b0) I8BE101CBEF6D2810BAC0C6F6AC8DA3B8 ; else if (IC79EC9A9F373F4B71374BDF6EDD31DE6
== 1'b1) I8BE101CBEF6D2810BAC0C6F6AC8DA3B8 ; else begin  if (I3DAC0A14B4001DD3A76D99313964C3AA ) I10F60E589450CD09FF7A498641DE26F8
<= {IB7D40CABAAA60621C763075C02B43B42 {1'b0}}; else begin if (I6316F5248B07D9065FBC7D67EDADC4EE ) I10F60E589450CD09FF7A498641DE26F8
<= (I10F60E589450CD09FF7A498641DE26F8 == (ID4C318F5AC8B6BE2D0E1091653FE0983 - 1)) ? {IB7D40CABAAA60621C763075C02B43B42 {1'b0}}
: (I10F60E589450CD09FF7A498641DE26F8 + 1); end  I102EDFAABB65014FC78C55AF4345F765 = {I6316F5248B07D9065FBC7D67EDADC4EE ,
I2FAC1854542B2B806297DF5B4733F9D2 }; case (I102EDFAABB65014FC78C55AF4345F765 ) 2'b01: begin I4FD65DDA0EDE2F39B09EF91789B31572
<= (IDDFF27981262750D43304A01A2EBF659 >= I1AF585FFD3730CB75D8EA561C736B279 ) ? 1'b0 : I4FD65DDA0EDE2F39B09EF91789B31572 ;
IDDFF27981262750D43304A01A2EBF659 <= IDDFF27981262750D43304A01A2EBF659 + ID4C318F5AC8B6BE2D0E1091653FE0983 ; I00CE0BA4F77A2426865D797055E4C98A
<= 1'b0; ID312B626B7C881C1A5210FC08BB95856 <= (I5C6C6CD7723900C21B3A76E887CEE164 == I64BB723AC8F87F7AEBA73BF190ED5F8F )
? I00CE0BA4F77A2426865D797055E4C98A : 1'b0; end 2'b10: begin I4FD65DDA0EDE2F39B09EF91789B31572 <= (IDDFF27981262750D43304A01A2EBF659
== IB011AB9176BFCCD54AFA433401B9CC28 ) ? 1'b1 : I4FD65DDA0EDE2F39B09EF91789B31572 ; IDDFF27981262750D43304A01A2EBF659
<= IDDFF27981262750D43304A01A2EBF659 - 1; I00CE0BA4F77A2426865D797055E4C98A <= I00CE0BA4F77A2426865D797055E4C98A
| ((IDDFF27981262750D43304A01A2EBF659 == 1) ? 1'b1 : 1'b0); ID312B626B7C881C1A5210FC08BB95856 <= (IDDFF27981262750D43304A01A2EBF659
== 2) ? 1'b1 : 1'b0; end 2'b11: begin I4FD65DDA0EDE2F39B09EF91789B31572 <= (IDDFF27981262750D43304A01A2EBF659 >=
I1AF585FFD3730CB75D8EA561C736B279 ) ? 1'b0 : I4FD65DDA0EDE2F39B09EF91789B31572 ; IDDFF27981262750D43304A01A2EBF659
<= IDDFF27981262750D43304A01A2EBF659 + (ID4C318F5AC8B6BE2D0E1091653FE0983 - 1); I00CE0BA4F77A2426865D797055E4C98A
<= 1'b0; ID312B626B7C881C1A5210FC08BB95856 <= (ID4C318F5AC8B6BE2D0E1091653FE0983 == 2) ? I00CE0BA4F77A2426865D797055E4C98A
: 1'b0; end endcase  ICA80E74165E79AFA565A1A052BE49F09 = {I38F39AED09C0507E780D3D35EA7FA06B , I2FAC1854542B2B806297DF5B4733F9D2 };
case (ICA80E74165E79AFA565A1A052BE49F09 ) 2'b01: begin I01F907CE74154BFFA0C1437099B21186 <= (IE1A203A1BCBBA5F947F638C3DFB65BF8
== I41D54753579217A07881641483914F62 ) ? 1'b1 : I01F907CE74154BFFA0C1437099B21186 ; ID079750A1760FEED5898B26A23289BAD
<= ID079750A1760FEED5898B26A23289BAD | ((IE1A203A1BCBBA5F947F638C3DFB65BF8 == 1) ? 1'b1 : 1'b0); IE1A203A1BCBBA5F947F638C3DFB65BF8
<= IE1A203A1BCBBA5F947F638C3DFB65BF8 - 1; I28ACD74043EE392893ABFA4360DDCD11 <= (IE1A203A1BCBBA5F947F638C3DFB65BF8
== 2) ? 1'b1 : 1'b0; end 2'b10: begin I01F907CE74154BFFA0C1437099B21186 <= (IE1A203A1BCBBA5F947F638C3DFB65BF8 ==
IC123CC1DD854BDF232C22DA342143DED ) ? 1'b0 : I01F907CE74154BFFA0C1437099B21186 ; ID079750A1760FEED5898B26A23289BAD
<= 1'b0; IE1A203A1BCBBA5F947F638C3DFB65BF8 <= IE1A203A1BCBBA5F947F638C3DFB65BF8 + 1; I28ACD74043EE392893ABFA4360DDCD11
<= ID079750A1760FEED5898B26A23289BAD ; end endcase    I69053399285CDFC39ECE32CB2CD079E5 = {I61018042B0489325A4CD993FF565603E ,
I6316F5248B07D9065FBC7D67EDADC4EE }; case (I69053399285CDFC39ECE32CB2CD079E5 ) 2'b01 : begin IDDCC249EE71726DC9EB38B3A433C91DB
<= IDDCC249EE71726DC9EB38B3A433C91DB - 1; I08DEC2092892554154AF13365E22F12A <= I08DEC2092892554154AF13365E22F12A
| ((IDDCC249EE71726DC9EB38B3A433C91DB == 1) ? 1'b1 : 1'b0); I6BE22F51BE43138B31F588DD2D062E1F <= 1'b0; end 2'b10
: begin IDDCC249EE71726DC9EB38B3A433C91DB <= IDDCC249EE71726DC9EB38B3A433C91DB + 1; I08DEC2092892554154AF13365E22F12A
<= 1'b0; I6BE22F51BE43138B31F588DD2D062E1F <= I6BE22F51BE43138B31F588DD2D062E1F | ((IDDCC249EE71726DC9EB38B3A433C91DB
== (I61D0345D311EC6FFC08DDDECE5F6127A - 1)) ? 1'b1 : 1'b0); end endcase  I07E46217B3640C9CD06BF9B9D5D78F68 <= I169F661B2921E0FA4AFB7C3794399862 ;
I7A2B537BEB4654059703B476744C6D18 <= I87FD0B6E6C89D593796D3B1F631D5100 ; I169F661B2921E0FA4AFB7C3794399862 <= I38F39AED09C0507E780D3D35EA7FA06B ;
I87FD0B6E6C89D593796D3B1F631D5100 <= I6316F5248B07D9065FBC7D67EDADC4EE ; I2E321486CBD81F71439B76F5D5BDCD93 <= I07E46217B3640C9CD06BF9B9D5D78F68
| I7A2B537BEB4654059703B476744C6D18 ; if (I38F39AED09C0507E780D3D35EA7FA06B == 1'b1) I3283453B42BD77672B8ACE724ACDA314
<= I3283453B42BD77672B8ACE724ACDA314 + 1; if (I2FAC1854542B2B806297DF5B4733F9D2 == 1'b1) IF8FA22381AE98928C01C1A8EF2CB0DC6
<= IF8FA22381AE98928C01C1A8EF2CB0DC6 + 1; if (I07E46217B3640C9CD06BF9B9D5D78F68 ) I134B7C80786213E899F61495BA54C91C
<= I1A61D2CA45ECC28270C28826CD87FEC3 ; else begin if (I7A2B537BEB4654059703B476744C6D18 ) I134B7C80786213E899F61495BA54C91C [I5C6C6CD7723900C21B3A76E887CEE164
- 1:0] <= I134B7C80786213E899F61495BA54C91C [I5C6C6CD7723900C21B3A76E887CEE164 - 1:0] >> I64BB723AC8F87F7AEBA73BF190ED5F8F ;
end end  end  end  endgenerate endmodule 
  module I2AA06444A0CB39074E17E74C913F2C98 # (parameter I7292F55C07BFD7FB8A60D29FFC186275 = 32, parameter I61D0345D311EC6FFC08DDDECE5F6127A
= 256 ) ( input wire ICCFB0F435B37370076102F325BC08D20 , input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire
IC79EC9A9F373F4B71374BDF6EDD31DE6 , input wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] ICFCA96AB1A120108CD0A9879E0F76EA8 ,
input wire ID8853B025150C80EE45BBA98E5BEA3A8 , input wire IF74C86FAF44E1757FDA146FCB1E10641 , input wire IA35D59E2E0D340C8C3D5ADB905E70579 ,
output wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] I125028C7446331521D0434C10E8B0007 , output wire I0D04F33C419DDB2EC0886F4409AB9A96 ,
output wire I585F74DE05DD9C1C7070D6B4F6E181C2 );  localparam I129D9485097D939AE1EF75F276EE6777 = 3; localparam IA14D7EA1BC849EB02A3E3D303AB9B071
= $clog2(I129D9485097D939AE1EF75F276EE6777 + 1); localparam I2F8DC10449A1F24468235753BBC3B988 = $clog2(I61D0345D311EC6FFC08DDDECE5F6127A
+ 1); localparam IF35F7B506981B2912E2486B227CB8871 = I7292F55C07BFD7FB8A60D29FFC186275 ;  reg [IF35F7B506981B2912E2486B227CB8871
- 1:0] I1140D78382474719F5279279A4E83ED5 [I129D9485097D939AE1EF75F276EE6777 - 1:0]; reg [I2F8DC10449A1F24468235753BBC3B988
- 1:0] I5206E2A6DE63CEC269DA56EACEB56A16 ; reg [IA14D7EA1BC849EB02A3E3D303AB9B071 - 1:0] IC6479B27A88B8B2D8B534765698B00EE ;
wire IF344AC55B7250509D3E5EC9317D747A5 ; wire I367E5D13940F83603F2CC8084CDC75AC ; wire I8873306A816AEB7F68F343867D02E5B8 ;
 assign I125028C7446331521D0434C10E8B0007 = (IC6479B27A88B8B2D8B534765698B00EE ) ? I1140D78382474719F5279279A4E83ED5 [IC6479B27A88B8B2D8B534765698B00EE
- 1] : ICFCA96AB1A120108CD0A9879E0F76EA8 ; assign I0D04F33C419DDB2EC0886F4409AB9A96 = I8873306A816AEB7F68F343867D02E5B8 ;
assign I585F74DE05DD9C1C7070D6B4F6E181C2 = (IC6479B27A88B8B2D8B534765698B00EE ) ? ~IF74C86FAF44E1757FDA146FCB1E10641
: IA35D59E2E0D340C8C3D5ADB905E70579 ;  assign IF344AC55B7250509D3E5EC9317D747A5 = (IC6479B27A88B8B2D8B534765698B00EE )
? ~IF74C86FAF44E1757FDA146FCB1E10641 : 1'b0; assign I367E5D13940F83603F2CC8084CDC75AC = (IF74C86FAF44E1757FDA146FCB1E10641
& IA35D59E2E0D340C8C3D5ADB905E70579 ) | (IF344AC55B7250509D3E5EC9317D747A5 & IA35D59E2E0D340C8C3D5ADB905E70579 );
assign I8873306A816AEB7F68F343867D02E5B8 = (IF74C86FAF44E1757FDA146FCB1E10641 ) ? 1'b0 : (ID8853B025150C80EE45BBA98E5BEA3A8
| (|I5206E2A6DE63CEC269DA56EACEB56A16 ));  generate if (1'b1) begin : I8CDDE92DE2910086C77F2B20C50D61C7 reg [1:0]
I151EFB3B054C018111728D0669873D94 ; reg [1:0] I7B20D86E7F1979C68D189FA6BA2F30A2 ; integer IC12312890F81D79D8CED15EE1E99727F ;
always @(posedge ICCFB0F435B37370076102F325BC08D20 or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin if (I9ED2A9117D3AEAF54CBA7AD69083BCB7
== 1'b0) begin I5206E2A6DE63CEC269DA56EACEB56A16 <= {I2F8DC10449A1F24468235753BBC3B988 {1'b0}}; IC6479B27A88B8B2D8B534765698B00EE
<= {IA14D7EA1BC849EB02A3E3D303AB9B071 {1'b0}}; for (IC12312890F81D79D8CED15EE1E99727F = 0; IC12312890F81D79D8CED15EE1E99727F
< I129D9485097D939AE1EF75F276EE6777 ; IC12312890F81D79D8CED15EE1E99727F = IC12312890F81D79D8CED15EE1E99727F + 1)
I1140D78382474719F5279279A4E83ED5 [IC12312890F81D79D8CED15EE1E99727F ] <= {IF35F7B506981B2912E2486B227CB8871 {1'b0}};
end else if (IC79EC9A9F373F4B71374BDF6EDD31DE6 == 1'b1) begin I5206E2A6DE63CEC269DA56EACEB56A16 <= {I2F8DC10449A1F24468235753BBC3B988 {1'b0}};
IC6479B27A88B8B2D8B534765698B00EE <= {IA14D7EA1BC849EB02A3E3D303AB9B071 {1'b0}}; for (IC12312890F81D79D8CED15EE1E99727F
= 0; IC12312890F81D79D8CED15EE1E99727F < I129D9485097D939AE1EF75F276EE6777 ; IC12312890F81D79D8CED15EE1E99727F =
IC12312890F81D79D8CED15EE1E99727F + 1) I1140D78382474719F5279279A4E83ED5 [IC12312890F81D79D8CED15EE1E99727F ] <=
{IF35F7B506981B2912E2486B227CB8871 {1'b0}}; end else begin  I7B20D86E7F1979C68D189FA6BA2F30A2 = {IF74C86FAF44E1757FDA146FCB1E10641 ,
ID8853B025150C80EE45BBA98E5BEA3A8 }; case (I7B20D86E7F1979C68D189FA6BA2F30A2 ) 2'b00 : begin I5206E2A6DE63CEC269DA56EACEB56A16
<= (I5206E2A6DE63CEC269DA56EACEB56A16 == 0) ? I5206E2A6DE63CEC269DA56EACEB56A16 : I5206E2A6DE63CEC269DA56EACEB56A16
- 1; end 2'b11 : begin I5206E2A6DE63CEC269DA56EACEB56A16 <= (I5206E2A6DE63CEC269DA56EACEB56A16 == I61D0345D311EC6FFC08DDDECE5F6127A )
? I5206E2A6DE63CEC269DA56EACEB56A16 : I5206E2A6DE63CEC269DA56EACEB56A16 + 1; end endcase  I151EFB3B054C018111728D0669873D94
= {IF344AC55B7250509D3E5EC9317D747A5 , I367E5D13940F83603F2CC8084CDC75AC }; case (I151EFB3B054C018111728D0669873D94 )
2'b01 : begin I1140D78382474719F5279279A4E83ED5 [0] <= ICFCA96AB1A120108CD0A9879E0F76EA8 ; IC6479B27A88B8B2D8B534765698B00EE
<= (IC6479B27A88B8B2D8B534765698B00EE == I129D9485097D939AE1EF75F276EE6777 ) ? IC6479B27A88B8B2D8B534765698B00EE
: IC6479B27A88B8B2D8B534765698B00EE + 1; for (IC12312890F81D79D8CED15EE1E99727F = 1; IC12312890F81D79D8CED15EE1E99727F
< I129D9485097D939AE1EF75F276EE6777 ; IC12312890F81D79D8CED15EE1E99727F = IC12312890F81D79D8CED15EE1E99727F + 1)
I1140D78382474719F5279279A4E83ED5 [IC12312890F81D79D8CED15EE1E99727F ] <= I1140D78382474719F5279279A4E83ED5 [IC12312890F81D79D8CED15EE1E99727F
- 1]; end 2'b10 : begin IC6479B27A88B8B2D8B534765698B00EE <= (IC6479B27A88B8B2D8B534765698B00EE ) ? IC6479B27A88B8B2D8B534765698B00EE
- 1 : 0; end 2'b11 : begin I1140D78382474719F5279279A4E83ED5 [0] <= ICFCA96AB1A120108CD0A9879E0F76EA8 ; for (IC12312890F81D79D8CED15EE1E99727F
= 1; IC12312890F81D79D8CED15EE1E99727F < I129D9485097D939AE1EF75F276EE6777 ; IC12312890F81D79D8CED15EE1E99727F =
IC12312890F81D79D8CED15EE1E99727F + 1) I1140D78382474719F5279279A4E83ED5 [IC12312890F81D79D8CED15EE1E99727F ] <=
I1140D78382474719F5279279A4E83ED5 [IC12312890F81D79D8CED15EE1E99727F - 1]; end endcase end end  end  endgenerate
endmodule
 `timescale 1 ns / 1 ps
module IF50ADBFC5F4E76B680AD98E97599279A # (parameter I424986699EB154C420BDB6FB59A8DA77 = 4, parameter I5D7F61632782AFE440ADE65900D53412
= 4, parameter I61D0345D311EC6FFC08DDDECE5F6127A = 256 ) ( input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input
wire ICCFB0F435B37370076102F325BC08D20 , input wire IC79EC9A9F373F4B71374BDF6EDD31DE6 , input wire ID8853B025150C80EE45BBA98E5BEA3A8 ,
input wire I22B24791BA0E7AA2C686B1B2D776C636 , output wire [$clog2(I61D0345D311EC6FFC08DDDECE5F6127A ) - 1:0] I79D313D86841E5141E7629EA606D7AE9 ,
output wire I11CEFC90537A67CD1FF01400245362F2 , output wire [$clog2(I61D0345D311EC6FFC08DDDECE5F6127A + 1) - 1:0]
ID7FCE45A65ADDB17F91F73A1B506BB5B , output wire I8BB939FF2AFDE7B2A1E480DCB61CE354 , output wire I41C63F948E534C7ED9F2471A44C922B2 ,
output wire I585F74DE05DD9C1C7070D6B4F6E181C2 , output wire [$clog2(I61D0345D311EC6FFC08DDDECE5F6127A ) - 1:0] I38B1AC532E13E69B05492C67EC7070BB ,
output wire I705C64753A50CDA034B5ACB332D71768 , output wire [$clog2(I61D0345D311EC6FFC08DDDECE5F6127A + 1) - 1:0]
I233E0C0C8E5150F0CD8258F276D93942 , output wire I102322A55721851004CB8E1F6AB50BDE , output wire IBE0D6810EBD63B5C428623C578CF6D3A ,
output wire I115E90220158F08B0465E99D7F2561D3 );  localparam I36A1B4EB5B5564A6ED7EA4D42856EFB4 = $clog2(I61D0345D311EC6FFC08DDDECE5F6127A );
localparam I2F8DC10449A1F24468235753BBC3B988 = $clog2(I61D0345D311EC6FFC08DDDECE5F6127A + 1); localparam I1AF585FFD3730CB75D8EA561C736B279
= I424986699EB154C420BDB6FB59A8DA77 ; localparam IB011AB9176BFCCD54AFA433401B9CC28 = I424986699EB154C420BDB6FB59A8DA77
+ 1; localparam IC123CC1DD854BDF232C22DA342143DED = I5D7F61632782AFE440ADE65900D53412 ; localparam I41D54753579217A07881641483914F62
= I5D7F61632782AFE440ADE65900D53412 + 1;  reg [I36A1B4EB5B5564A6ED7EA4D42856EFB4 - 1:0] I3283453B42BD77672B8ACE724ACDA314 ;
reg [I36A1B4EB5B5564A6ED7EA4D42856EFB4 - 1:0] IF8FA22381AE98928C01C1A8EF2CB0DC6 ; reg I68525D8B661ABC93EC5BB1B92FE9724E ;
reg I4FD65DDA0EDE2F39B09EF91789B31572 ; reg [I2F8DC10449A1F24468235753BBC3B988 - 1:0] IDDFF27981262750D43304A01A2EBF659 ;
reg I00CE0BA4F77A2426865D797055E4C98A ; reg ID312B626B7C881C1A5210FC08BB95856 ; reg [I2F8DC10449A1F24468235753BBC3B988
- 1:0] I150212E44B1214E167CE3FB321CC3459 ; reg I05305DB38B053FE192F0B71598347D85 ; reg I01F907CE74154BFFA0C1437099B21186 ;
reg [I2F8DC10449A1F24468235753BBC3B988 - 1:0] IE1A203A1BCBBA5F947F638C3DFB65BF8 ; reg ID079750A1760FEED5898B26A23289BAD ;
reg I28ACD74043EE392893ABFA4360DDCD11 ; wire I2C3263714ADF8DC5044612F1D1CA7C60 ; wire I0F5257612C50B0E646400AEA2A64E768 ;
wire I2FAC1854542B2B806297DF5B4733F9D2 ;  assign I79D313D86841E5141E7629EA606D7AE9 = I3283453B42BD77672B8ACE724ACDA314 ;
assign I11CEFC90537A67CD1FF01400245362F2 = I4FD65DDA0EDE2F39B09EF91789B31572 ; assign ID7FCE45A65ADDB17F91F73A1B506BB5B
= IDDFF27981262750D43304A01A2EBF659 ; assign I8BB939FF2AFDE7B2A1E480DCB61CE354 = I00CE0BA4F77A2426865D797055E4C98A ;
assign I41C63F948E534C7ED9F2471A44C922B2 = ID312B626B7C881C1A5210FC08BB95856 ; assign I585F74DE05DD9C1C7070D6B4F6E181C2
= I05305DB38B053FE192F0B71598347D85 ; assign I38B1AC532E13E69B05492C67EC7070BB = IF8FA22381AE98928C01C1A8EF2CB0DC6 ;
assign I705C64753A50CDA034B5ACB332D71768 = I01F907CE74154BFFA0C1437099B21186 ; assign I233E0C0C8E5150F0CD8258F276D93942
= IE1A203A1BCBBA5F947F638C3DFB65BF8 ; assign I102322A55721851004CB8E1F6AB50BDE = I2FAC1854542B2B806297DF5B4733F9D2 ;
assign IBE0D6810EBD63B5C428623C578CF6D3A = ID079750A1760FEED5898B26A23289BAD ; assign I115E90220158F08B0465E99D7F2561D3
= I28ACD74043EE392893ABFA4360DDCD11 ;  assign I2C3263714ADF8DC5044612F1D1CA7C60 = ID8853B025150C80EE45BBA98E5BEA3A8
& ~I00CE0BA4F77A2426865D797055E4C98A ; assign I0F5257612C50B0E646400AEA2A64E768 = (I150212E44B1214E167CE3FB321CC3459
> 0) ? 1'b1 : 1'b0; assign I2FAC1854542B2B806297DF5B4733F9D2 = I22B24791BA0E7AA2C686B1B2D776C636 & ~ID079750A1760FEED5898B26A23289BAD ;
 generate if (1'b1) begin : I8CDDE92DE2910086C77F2B20C50D61C7 reg [1:0] I151EFB3B054C018111728D0669873D94 ; reg
[1:0] I102EDFAABB65014FC78C55AF4345F765 ; reg [1:0] I69053399285CDFC39ECE32CB2CD079E5 ; reg [1:0] ICA80E74165E79AFA565A1A052BE49F09 ;
integer IC12312890F81D79D8CED15EE1E99727F ; task I8BE101CBEF6D2810BAC0C6F6AC8DA3B8 ; begin I3283453B42BD77672B8ACE724ACDA314
<= 0; IF8FA22381AE98928C01C1A8EF2CB0DC6 <= 0; I68525D8B661ABC93EC5BB1B92FE9724E <= 1'b0; I4FD65DDA0EDE2F39B09EF91789B31572
<= 1'b0; I00CE0BA4F77A2426865D797055E4C98A <= 1'b1; IDDFF27981262750D43304A01A2EBF659 <= 0; ID312B626B7C881C1A5210FC08BB95856
<= 1'b0; I150212E44B1214E167CE3FB321CC3459 <= 0; I05305DB38B053FE192F0B71598347D85 <= 1'b0; I01F907CE74154BFFA0C1437099B21186
<= 1'b0; ID079750A1760FEED5898B26A23289BAD <= 1'b0; IE1A203A1BCBBA5F947F638C3DFB65BF8 <= I61D0345D311EC6FFC08DDDECE5F6127A ;
I28ACD74043EE392893ABFA4360DDCD11 <= 1'b0; end endtask always @(posedge ICCFB0F435B37370076102F325BC08D20 or negedge
I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin if (I9ED2A9117D3AEAF54CBA7AD69083BCB7 == 1'b0) I8BE101CBEF6D2810BAC0C6F6AC8DA3B8 ;
else if (IC79EC9A9F373F4B71374BDF6EDD31DE6 == 1'b1) I8BE101CBEF6D2810BAC0C6F6AC8DA3B8 ; else begin I102EDFAABB65014FC78C55AF4345F765
= {I2C3263714ADF8DC5044612F1D1CA7C60 , I2FAC1854542B2B806297DF5B4733F9D2 }; case (I102EDFAABB65014FC78C55AF4345F765 )
2'b01: begin I4FD65DDA0EDE2F39B09EF91789B31572 <= (IDDFF27981262750D43304A01A2EBF659 == I1AF585FFD3730CB75D8EA561C736B279 )
? 1'b0 : I4FD65DDA0EDE2F39B09EF91789B31572 ; I00CE0BA4F77A2426865D797055E4C98A <= 1'b0; IDDFF27981262750D43304A01A2EBF659
<= IDDFF27981262750D43304A01A2EBF659 + 1; ID312B626B7C881C1A5210FC08BB95856 <= I00CE0BA4F77A2426865D797055E4C98A ;
end 2'b10: begin I4FD65DDA0EDE2F39B09EF91789B31572 <= (IDDFF27981262750D43304A01A2EBF659 == IB011AB9176BFCCD54AFA433401B9CC28 )
? 1'b1 : I4FD65DDA0EDE2F39B09EF91789B31572 ; I00CE0BA4F77A2426865D797055E4C98A <= I00CE0BA4F77A2426865D797055E4C98A
| ((IDDFF27981262750D43304A01A2EBF659 == 1) ? 1'b1 : 1'b0); IDDFF27981262750D43304A01A2EBF659 <= IDDFF27981262750D43304A01A2EBF659
- 1; ID312B626B7C881C1A5210FC08BB95856 <= (IDDFF27981262750D43304A01A2EBF659 == 2) ? 1'b1 : 1'b0; end endcase  ICA80E74165E79AFA565A1A052BE49F09
= {I2C3263714ADF8DC5044612F1D1CA7C60 , I2FAC1854542B2B806297DF5B4733F9D2 }; case (ICA80E74165E79AFA565A1A052BE49F09 )
2'b01: begin I01F907CE74154BFFA0C1437099B21186 <= (IE1A203A1BCBBA5F947F638C3DFB65BF8 == I41D54753579217A07881641483914F62 )
? 1'b1 : I01F907CE74154BFFA0C1437099B21186 ; ID079750A1760FEED5898B26A23289BAD <= ID079750A1760FEED5898B26A23289BAD
| ((IE1A203A1BCBBA5F947F638C3DFB65BF8 == 1) ? 1'b1 : 1'b0); IE1A203A1BCBBA5F947F638C3DFB65BF8 <= IE1A203A1BCBBA5F947F638C3DFB65BF8
- 1; I28ACD74043EE392893ABFA4360DDCD11 <= (IE1A203A1BCBBA5F947F638C3DFB65BF8 == 2) ? 1'b1 : 1'b0; end 2'b10: begin
I01F907CE74154BFFA0C1437099B21186 <= (IE1A203A1BCBBA5F947F638C3DFB65BF8 == IC123CC1DD854BDF232C22DA342143DED ) ?
1'b0 : I01F907CE74154BFFA0C1437099B21186 ; ID079750A1760FEED5898B26A23289BAD <= 1'b0; IE1A203A1BCBBA5F947F638C3DFB65BF8
<= IE1A203A1BCBBA5F947F638C3DFB65BF8 + 1; I28ACD74043EE392893ABFA4360DDCD11 <= ID079750A1760FEED5898B26A23289BAD ;
end endcase   I69053399285CDFC39ECE32CB2CD079E5 = {I2C3263714ADF8DC5044612F1D1CA7C60 , I0F5257612C50B0E646400AEA2A64E768 };
case (I69053399285CDFC39ECE32CB2CD079E5 ) 2'b01 : begin I150212E44B1214E167CE3FB321CC3459 <= I150212E44B1214E167CE3FB321CC3459
- 1; end 2'b10 : begin I150212E44B1214E167CE3FB321CC3459 <= I150212E44B1214E167CE3FB321CC3459 + 1; end endcase 
I68525D8B661ABC93EC5BB1B92FE9724E <= I0F5257612C50B0E646400AEA2A64E768 ; I05305DB38B053FE192F0B71598347D85 <= I68525D8B661ABC93EC5BB1B92FE9724E ;
if (I0F5257612C50B0E646400AEA2A64E768 ) I3283453B42BD77672B8ACE724ACDA314 <= I3283453B42BD77672B8ACE724ACDA314 +
1; if (I2FAC1854542B2B806297DF5B4733F9D2 == 1'b1) IF8FA22381AE98928C01C1A8EF2CB0DC6 <= IF8FA22381AE98928C01C1A8EF2CB0DC6
+ 1; end  end  end  endgenerate endmodule 
  `timescale 1 ns / 1 ps 
module IF4FD65273243DC47A72869EEEA639DCD # (parameter I7292F55C07BFD7FB8A60D29FFC186275 = 32, parameter IB71844FFA3AB85FEF45EAB4D35395752
= 512, parameter I424986699EB154C420BDB6FB59A8DA77 = 4, parameter I5D7F61632782AFE440ADE65900D53412 = 4, parameter
I66C185998F46A7148163982E39BCD296 = "ecp3" ) ( input wire ICCFB0F435B37370076102F325BC08D20 , input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 ,
input wire IC79EC9A9F373F4B71374BDF6EDD31DE6 , input wire I48D61F5A0B5732A58912433B42CD9D0C , input wire [I7292F55C07BFD7FB8A60D29FFC186275
- 1:0] I04BC24D2B6403E54A64DE9E6C9ABAA2B , input wire IE315CDCA06C9620D5C0AB966E553F0C3 , output wire I11CEFC90537A67CD1FF01400245362F2 ,
output wire [$clog2(IB71844FFA3AB85FEF45EAB4D35395752 + 1) - 1:0] ID7FCE45A65ADDB17F91F73A1B506BB5B , output wire
[I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] I125028C7446331521D0434C10E8B0007 , output wire I8BB939FF2AFDE7B2A1E480DCB61CE354 ,
output wire I41C63F948E534C7ED9F2471A44C922B2 , output wire I585F74DE05DD9C1C7070D6B4F6E181C2 , output wire I705C64753A50CDA034B5ACB332D71768 ,
output wire [$clog2(IB71844FFA3AB85FEF45EAB4D35395752 + 1) - 1:0] I233E0C0C8E5150F0CD8258F276D93942 , output wire
IBE0D6810EBD63B5C428623C578CF6D3A , output wire I115E90220158F08B0465E99D7F2561D3 );  localparam integer I36A1B4EB5B5564A6ED7EA4D42856EFB4
= $clog2(IB71844FFA3AB85FEF45EAB4D35395752 ); localparam integer I2F8DC10449A1F24468235753BBC3B988 = $clog2(IB71844FFA3AB85FEF45EAB4D35395752
+ 1); localparam integer IF35F7B506981B2912E2486B227CB8871 = I7292F55C07BFD7FB8A60D29FFC186275 ;  wire [I36A1B4EB5B5564A6ED7EA4D42856EFB4
- 1:0] IC2A6ECC367E2C82B97E73A57A8A79E1A ; wire IF6E67DBB7CD3AAE309AE42CCEEB33046 ; wire [I2F8DC10449A1F24468235753BBC3B988
- 1:0] I366D7D477BCE878309C2A4C6F4920631 ; wire I60B15FF62AA99717C8B7DA7D6912D281 ; wire ICB86B570A185B89048AE76A09444BA41 ;
wire IA6BBDC90BCC6EF2E35BFA8D709343BF3 ; wire [I36A1B4EB5B5564A6ED7EA4D42856EFB4 - 1:0] I5631F39935597168A2C9D3656C66CB5C ;
wire I0E620501249C5CFBF447631D04D33715 ; wire [I2F8DC10449A1F24468235753BBC3B988 - 1:0] I1E2790529716BDA31237F724D6F3C1DA ;
wire I25891FD4BF8EA7F9051CE324A21ED31E ; wire I366EB0B781FD462E1BDC374519E76C20 ; wire IF63FD497AC79A293EAC51C0F982F9AD3 ;
wire [IF35F7B506981B2912E2486B227CB8871 - 1:0] I2CA1A324143051A0AFDEFB54659C657C ; wire I4AE98FF3DA4D5A5EE68F8A14D9D781F4 ;
 assign I11CEFC90537A67CD1FF01400245362F2 = IF6E67DBB7CD3AAE309AE42CCEEB33046 ; assign ID7FCE45A65ADDB17F91F73A1B506BB5B
= I366D7D477BCE878309C2A4C6F4920631 ; assign I125028C7446331521D0434C10E8B0007 = I2CA1A324143051A0AFDEFB54659C657C ;
assign I8BB939FF2AFDE7B2A1E480DCB61CE354 = I60B15FF62AA99717C8B7DA7D6912D281 ; assign I41C63F948E534C7ED9F2471A44C922B2
= ICB86B570A185B89048AE76A09444BA41 ; assign I585F74DE05DD9C1C7070D6B4F6E181C2 = IA6BBDC90BCC6EF2E35BFA8D709343BF3 ;
assign I705C64753A50CDA034B5ACB332D71768 = I0E620501249C5CFBF447631D04D33715 ; assign I233E0C0C8E5150F0CD8258F276D93942
= I1E2790529716BDA31237F724D6F3C1DA ; assign IBE0D6810EBD63B5C428623C578CF6D3A = I366EB0B781FD462E1BDC374519E76C20 ;
assign I115E90220158F08B0465E99D7F2561D3 = IF63FD497AC79A293EAC51C0F982F9AD3 ;  assign I4AE98FF3DA4D5A5EE68F8A14D9D781F4
= ~I9ED2A9117D3AEAF54CBA7AD69083BCB7 ;  IF50ADBFC5F4E76B680AD98E97599279A #( .I424986699EB154C420BDB6FB59A8DA77
(I424986699EB154C420BDB6FB59A8DA77 ), .I5D7F61632782AFE440ADE65900D53412 (I5D7F61632782AFE440ADE65900D53412 ), .I61D0345D311EC6FFC08DDDECE5F6127A
(IB71844FFA3AB85FEF45EAB4D35395752 ) ) IB420C4D1279F971E867FA537CA4D6E82 ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ),
.I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .IC79EC9A9F373F4B71374BDF6EDD31DE6 (IC79EC9A9F373F4B71374BDF6EDD31DE6 ),
.ID8853B025150C80EE45BBA98E5BEA3A8 (I48D61F5A0B5732A58912433B42CD9D0C ), .I22B24791BA0E7AA2C686B1B2D776C636 (IE315CDCA06C9620D5C0AB966E553F0C3 ),
.I79D313D86841E5141E7629EA606D7AE9 (IC2A6ECC367E2C82B97E73A57A8A79E1A ), .I11CEFC90537A67CD1FF01400245362F2 (IF6E67DBB7CD3AAE309AE42CCEEB33046 ),
.ID7FCE45A65ADDB17F91F73A1B506BB5B (I366D7D477BCE878309C2A4C6F4920631 ), .I8BB939FF2AFDE7B2A1E480DCB61CE354 (I60B15FF62AA99717C8B7DA7D6912D281 ),
.I41C63F948E534C7ED9F2471A44C922B2 (ICB86B570A185B89048AE76A09444BA41 ), .I585F74DE05DD9C1C7070D6B4F6E181C2 (IA6BBDC90BCC6EF2E35BFA8D709343BF3 ),
.I38B1AC532E13E69B05492C67EC7070BB (I5631F39935597168A2C9D3656C66CB5C ), .I705C64753A50CDA034B5ACB332D71768 (I0E620501249C5CFBF447631D04D33715 ),
.I102322A55721851004CB8E1F6AB50BDE (I25891FD4BF8EA7F9051CE324A21ED31E ), .I233E0C0C8E5150F0CD8258F276D93942 (I1E2790529716BDA31237F724D6F3C1DA ),
.IBE0D6810EBD63B5C428623C578CF6D3A (I366EB0B781FD462E1BDC374519E76C20 ), .I115E90220158F08B0465E99D7F2561D3 (IF63FD497AC79A293EAC51C0F982F9AD3 )
); pmi_ram_dp # ( .pmi_wr_addr_depth (IB71844FFA3AB85FEF45EAB4D35395752 ), .pmi_wr_addr_width (I36A1B4EB5B5564A6ED7EA4D42856EFB4 ),
.pmi_wr_data_width (IF35F7B506981B2912E2486B227CB8871 ), .pmi_rd_addr_depth (IB71844FFA3AB85FEF45EAB4D35395752 ),
.pmi_rd_addr_width (I36A1B4EB5B5564A6ED7EA4D42856EFB4 ), .pmi_rd_data_width (IF35F7B506981B2912E2486B227CB8871 ),
.pmi_regmode ("reg"), .pmi_family (I66C185998F46A7148163982E39BCD296 ), .module_type ("pmi_ram_dp") ) I32900CECD80193336B4F376406D5DFF6
( .Data (I04BC24D2B6403E54A64DE9E6C9ABAA2B ), .RdAddress (IC2A6ECC367E2C82B97E73A57A8A79E1A ), .RdClockEn (1'b1),
.RdClock (ICCFB0F435B37370076102F325BC08D20 ), .Reset (I4AE98FF3DA4D5A5EE68F8A14D9D781F4 ), .WE (I25891FD4BF8EA7F9051CE324A21ED31E ),
.WrAddress (I5631F39935597168A2C9D3656C66CB5C ), .WrClockEn (1'b1), .WrClock (ICCFB0F435B37370076102F325BC08D20 ),
.Q (I2CA1A324143051A0AFDEFB54659C657C ) ); endmodule 
  module I792C47F7E7D7705A2329EEB04CA92E91 ( input wire ICCFB0F435B37370076102F325BC08D20 , input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 ,
input wire I93AE636CE82DE94CB11ACCF59F8C2254 , input wire [15:0] I2AED852F071D7FF5A04BEFAF4E7F3B0F , input wire
I9B9FF20B523F68871F4D27848F9B4E44 , input wire I694FF88E6CB22CE905A2A9A9E00AF7F1 , output wire [31:0] IF249B786312150CAA567D0B3F1DC760E ,
output wire I99A7C01D853D4CD1BF86EA17B055AE82 , output wire IAB7D8322CEA20D7B2FC0EF19A061CB19 , output wire I14B85FB28FCEF458E6F9665F2960F9A2 ,
output wire [31:0] I528AB843F22B93013A3EAA53871813E4 , output wire I55EF6D8E66D2B56872BA18F8A67DBCC9 , output wire
ICF9485DAA5CD85FD9CF3AB9F6898D8FC , output wire I3E859D8CBD08E747693AC2BA98F2B947 ); `include "pcisig_constants.v"
 reg IE97C1EAB688C29EF293B3533128589AD ; reg I7E9F566F873687A02EB36D908875E0CE ; reg [2:0] I31B6AE50934C66C240CC08D3DC502236 ;
reg I9C1F19035765F165886CDE9ADA8857F3 ; reg I54BE80AB8C90F3E5819921EF5354732A ; reg IDA82F4C78A43B62E1C09ED19A1443221 ;
reg IB4FFC03833EA896621BFDB5DCC2E1B6D ; reg [15:0] IA9505001B62C5345479286119EE12C81 ; reg IE9F53C1FA095EA11A4F2438E8D110DCB ;
reg I91DDB59BA2C93482521ADEF2F41C8F5F ; reg [31:0] ID5AB6F130EBFA08B3BFFD3C140B232D7 ; reg I7CDEBB8EE6259E09FDB23A8CB9153F7B ;
reg I6DC757833BFBECB509EE1BB6128BCB2D ; reg I08158090CAF768A22FBFA7B602DA8EE9 ; reg I0935F33573E9008AC6C383C6271492EC ;
wire IE12D7FB0707DA0B72DA8BD64B6FAEFEB ;  assign IF249B786312150CAA567D0B3F1DC760E = {ID5AB6F130EBFA08B3BFFD3C140B232D7 [7:0],
ID5AB6F130EBFA08B3BFFD3C140B232D7 [15:8], ID5AB6F130EBFA08B3BFFD3C140B232D7 [23:16], ID5AB6F130EBFA08B3BFFD3C140B232D7 [31:24]};
assign I99A7C01D853D4CD1BF86EA17B055AE82 = I7E9F566F873687A02EB36D908875E0CE ; assign IAB7D8322CEA20D7B2FC0EF19A061CB19
= I31B6AE50934C66C240CC08D3DC502236 [2]; assign I14B85FB28FCEF458E6F9665F2960F9A2 = I9C1F19035765F165886CDE9ADA8857F3 ;
assign I528AB843F22B93013A3EAA53871813E4 = ID5AB6F130EBFA08B3BFFD3C140B232D7 ; assign I55EF6D8E66D2B56872BA18F8A67DBCC9
= I7CDEBB8EE6259E09FDB23A8CB9153F7B ; assign ICF9485DAA5CD85FD9CF3AB9F6898D8FC = I6DC757833BFBECB509EE1BB6128BCB2D ;
assign I3E859D8CBD08E747693AC2BA98F2B947 = I0935F33573E9008AC6C383C6271492EC ;  assign IE12D7FB0707DA0B72DA8BD64B6FAEFEB
= ((IA9505001B62C5345479286119EE12C81 [15:8] == I6A62FD6104E281B8714322DB8CCB5FE3 ) || (IA9505001B62C5345479286119EE12C81 [15:8]
== I85B0192F2AC4464C88E2C93352FE6696 ) || (IA9505001B62C5345479286119EE12C81 [15:8] == I78DDE5821936F928E302A8BA3C3138EE )
|| (IA9505001B62C5345479286119EE12C81 [15:8] == I41F249A62806D544C38454CA2D10750D )) ? 1'b1 : 1'b0;  always @(posedge
ICCFB0F435B37370076102F325BC08D20 or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) if (~I9ED2A9117D3AEAF54CBA7AD69083BCB7 )
begin IE97C1EAB688C29EF293B3533128589AD <= 1'b0; I7E9F566F873687A02EB36D908875E0CE <= 1'b0; I31B6AE50934C66C240CC08D3DC502236
<= 3'b0; I9C1F19035765F165886CDE9ADA8857F3 <= 1'b0; I54BE80AB8C90F3E5819921EF5354732A <= 1'b0; IDA82F4C78A43B62E1C09ED19A1443221
<= 1'b0; IB4FFC03833EA896621BFDB5DCC2E1B6D <= 1'b0; IA9505001B62C5345479286119EE12C81 <= 16'b0; IE9F53C1FA095EA11A4F2438E8D110DCB
<= 1'b0; I91DDB59BA2C93482521ADEF2F41C8F5F <= 1'b0; ID5AB6F130EBFA08B3BFFD3C140B232D7 <= 32'b0; I7CDEBB8EE6259E09FDB23A8CB9153F7B
<= 1'b0; I6DC757833BFBECB509EE1BB6128BCB2D <= 1'b0; I08158090CAF768A22FBFA7B602DA8EE9 <= 1'b0; I0935F33573E9008AC6C383C6271492EC
<= 1'b0; end else begin IE97C1EAB688C29EF293B3533128589AD <= IE97C1EAB688C29EF293B3533128589AD & ~IE9F53C1FA095EA11A4F2438E8D110DCB ;
I9C1F19035765F165886CDE9ADA8857F3 <= 1'b0; I54BE80AB8C90F3E5819921EF5354732A <= I93AE636CE82DE94CB11ACCF59F8C2254 ;
IA9505001B62C5345479286119EE12C81 <= I2AED852F071D7FF5A04BEFAF4E7F3B0F ; IE9F53C1FA095EA11A4F2438E8D110DCB <= I9B9FF20B523F68871F4D27848F9B4E44 ;
I91DDB59BA2C93482521ADEF2F41C8F5F <= I694FF88E6CB22CE905A2A9A9E00AF7F1 ; I08158090CAF768A22FBFA7B602DA8EE9 <= I08158090CAF768A22FBFA7B602DA8EE9
& ~IE9F53C1FA095EA11A4F2438E8D110DCB ; I0935F33573E9008AC6C383C6271492EC <= 1'b0; if (I91DDB59BA2C93482521ADEF2F41C8F5F
& I54BE80AB8C90F3E5819921EF5354732A ) begin IE97C1EAB688C29EF293B3533128589AD <= IE12D7FB0707DA0B72DA8BD64B6FAEFEB ;
I7E9F566F873687A02EB36D908875E0CE <= IE12D7FB0707DA0B72DA8BD64B6FAEFEB ; I31B6AE50934C66C240CC08D3DC502236 <= 3'b0;
IDA82F4C78A43B62E1C09ED19A1443221 <= IA9505001B62C5345479286119EE12C81 [14]; IB4FFC03833EA896621BFDB5DCC2E1B6D <=
1'b1; I7CDEBB8EE6259E09FDB23A8CB9153F7B <= 1'b0; I6DC757833BFBECB509EE1BB6128BCB2D <= 1'b1; I08158090CAF768A22FBFA7B602DA8EE9
<= ~IE12D7FB0707DA0B72DA8BD64B6FAEFEB ; ID5AB6F130EBFA08B3BFFD3C140B232D7 [31:16] <= IA9505001B62C5345479286119EE12C81 ;
end if (IE97C1EAB688C29EF293B3533128589AD | I08158090CAF768A22FBFA7B602DA8EE9 ) begin IB4FFC03833EA896621BFDB5DCC2E1B6D
<= ~IB4FFC03833EA896621BFDB5DCC2E1B6D ; I7CDEBB8EE6259E09FDB23A8CB9153F7B <= IE9F53C1FA095EA11A4F2438E8D110DCB ;
if (IB4FFC03833EA896621BFDB5DCC2E1B6D ) begin I9C1F19035765F165886CDE9ADA8857F3 <= IE97C1EAB688C29EF293B3533128589AD ;
ID5AB6F130EBFA08B3BFFD3C140B232D7 [15:0] <= IA9505001B62C5345479286119EE12C81 ; I0935F33573E9008AC6C383C6271492EC
<= I08158090CAF768A22FBFA7B602DA8EE9 ; end else begin I7E9F566F873687A02EB36D908875E0CE <= I7E9F566F873687A02EB36D908875E0CE
& ~I31B6AE50934C66C240CC08D3DC502236 [1]; I31B6AE50934C66C240CC08D3DC502236 <= {I31B6AE50934C66C240CC08D3DC502236 [1:0],
(IDA82F4C78A43B62E1C09ED19A1443221 & IE97C1EAB688C29EF293B3533128589AD )}; I9C1F19035765F165886CDE9ADA8857F3 <=
1'b0; ID5AB6F130EBFA08B3BFFD3C140B232D7 [31:16] <= IA9505001B62C5345479286119EE12C81 ; I6DC757833BFBECB509EE1BB6128BCB2D
<= 1'b0; I0935F33573E9008AC6C383C6271492EC <= 1'b0; end end end endmodule 
  module IB48580D48DC6311D8E12B4626CE243D8 ( input wire ICCFB0F435B37370076102F325BC08D20 , input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 ,
input wire I93AE636CE82DE94CB11ACCF59F8C2254 , input wire [63:0] I2AED852F071D7FF5A04BEFAF4E7F3B0F , input wire
I9B9FF20B523F68871F4D27848F9B4E44 , input wire I694FF88E6CB22CE905A2A9A9E00AF7F1 , output wire IA05976160EBA6DEFAAAA66970A81B32D ,
output wire [63:0] IF249B786312150CAA567D0B3F1DC760E , output wire ID7EB8E74BC37FDF7521CAA3A6410AD1C , output wire
I0DE0BA1FE7C719C02C2286C7BB4E82EC , output wire [2:0] I22CD4A94B7889ACD9A7D67943BC18F3B , output wire [10:0] I4F75D3BA09A515DCAD40830FB24835A7 ,
output wire I14B85FB28FCEF458E6F9665F2960F9A2 , output wire [63:0] I528AB843F22B93013A3EAA53871813E4 , output wire
I55EF6D8E66D2B56872BA18F8A67DBCC9 , output wire ICF9485DAA5CD85FD9CF3AB9F6898D8FC , output wire I6CE3395345F58F9D860AC549C8AF1473
); `include "pcisig_constants.v" 
 localparam IE13B4590716ED954FC344B681DC7BBA6 = 2;  reg I6B994CECB5A77B313B1493CB67891E99 ; reg [63:0] I109D319C018EB616621364D94266DBCD ;
reg IBABAB34D868FD2B2C7A88C42E97BBE11 ; reg I265478FD9C844733CCACAB4D3F6F7A3F ; reg [2:0] IECFDE780B7B9CC7363547C818E204EBB ;
reg [10:0] I1B52D4A8BF5D40A682398CBEA678902A ; reg I9C1F19035765F165886CDE9ADA8857F3 ; reg I54BE80AB8C90F3E5819921EF5354732A ;
reg I586C583482F0FD3AF11293684F55AD76 ; reg I57B81EC60D40AFFA64B92817187C45D7 ; reg I028038B8A4E4CB73C6DD88AF8C0C9F3E ;
reg [IE13B4590716ED954FC344B681DC7BBA6 - 1:0] I46B34B7B5B0375E4DD3F84053E6360B7 ; reg [2:0] I7D0FD152081CEE292550C7730CCA5F75 ;
reg [10:0] I64D52FE53B2984CB9C38CC7D9230077D ; reg [63:0] IA9505001B62C5345479286119EE12C81 [IE13B4590716ED954FC344B681DC7BBA6
- 1:0]; reg [IE13B4590716ED954FC344B681DC7BBA6 - 1:0] IE9F53C1FA095EA11A4F2438E8D110DCB ; reg [IE13B4590716ED954FC344B681DC7BBA6
- 1:0] I6EEF1710176D9017BF7C396C5C2DDAD6 ; reg [63:0] I72AC15FBC2C6EF14364CFFBBB83E3AC0 ; reg [63:0] IFAB2125DC13DFE796F8D4DDBDFC09F4A ;
reg I9F845E1C893E9E4563815DFDDDFF7E5B ; reg I674E1FE7EB5BC40955A2009618388E94 ; reg I2A6B381FD8829A5C8BD04107C91C9378 ;
reg IE68E826F0832B729C0DA0FA2B2697E2E ; reg I3A905796D2783CA2AD55AEB4DA75441A ; reg I1A378769CCB13A524F53158EF54CADD0 ;
reg I5E5A9B8E7ABF32287F37CE45D050FE5F ; reg I1407533F2D3FCAAA5E6EC4C54A09AEB5 ; reg IE8B637460BB6B1FB35EB926F2D20C02B ;
reg [63:0] ID5AB6F130EBFA08B3BFFD3C140B232D7 ; reg I2D1CB7F5C024D3CED1F017A4D3BC1F55 ; wire IDA82F4C78A43B62E1C09ED19A1443221 ;
wire IE12D7FB0707DA0B72DA8BD64B6FAEFEB ; wire I049E6CF82F9492802746D564E2B88117 ; wire I0515522FF1EFD23C59D28B8F6AB3A424 ;
 assign IA05976160EBA6DEFAAAA66970A81B32D = I6B994CECB5A77B313B1493CB67891E99 ; assign IF249B786312150CAA567D0B3F1DC760E
= I109D319C018EB616621364D94266DBCD ; assign ID7EB8E74BC37FDF7521CAA3A6410AD1C = IBABAB34D868FD2B2C7A88C42E97BBE11 ;
assign I0DE0BA1FE7C719C02C2286C7BB4E82EC = I265478FD9C844733CCACAB4D3F6F7A3F ; assign I22CD4A94B7889ACD9A7D67943BC18F3B
= IECFDE780B7B9CC7363547C818E204EBB ; assign I4F75D3BA09A515DCAD40830FB24835A7 = I1B52D4A8BF5D40A682398CBEA678902A ;
assign I14B85FB28FCEF458E6F9665F2960F9A2 = I9C1F19035765F165886CDE9ADA8857F3 ; assign I528AB843F22B93013A3EAA53871813E4
= {ID5AB6F130EBFA08B3BFFD3C140B232D7 [31:0], ID5AB6F130EBFA08B3BFFD3C140B232D7 [63:32]}; assign I55EF6D8E66D2B56872BA18F8A67DBCC9
= IE9F53C1FA095EA11A4F2438E8D110DCB [1]; assign ICF9485DAA5CD85FD9CF3AB9F6898D8FC = I6EEF1710176D9017BF7C396C5C2DDAD6 [1];
assign I6CE3395345F58F9D860AC549C8AF1473 = IE8B637460BB6B1FB35EB926F2D20C02B ;  assign IDA82F4C78A43B62E1C09ED19A1443221
= IA9505001B62C5345479286119EE12C81 [0][62]; assign IE12D7FB0707DA0B72DA8BD64B6FAEFEB = ((IA9505001B62C5345479286119EE12C81 [0][63:56]
== I6A62FD6104E281B8714322DB8CCB5FE3 ) || (IA9505001B62C5345479286119EE12C81 [0][63:56] == I85B0192F2AC4464C88E2C93352FE6696 )
|| (IA9505001B62C5345479286119EE12C81 [0][63:56] == I78DDE5821936F928E302A8BA3C3138EE ) || (IA9505001B62C5345479286119EE12C81 [0][63:56]
== I41F249A62806D544C38454CA2D10750D )) ? 1'b1 : 1'b0; assign I049E6CF82F9492802746D564E2B88117 = (I2D1CB7F5C024D3CED1F017A4D3BC1F55
== 1'b1) ? IE9F53C1FA095EA11A4F2438E8D110DCB [1] : IE9F53C1FA095EA11A4F2438E8D110DCB [0]; assign I0515522FF1EFD23C59D28B8F6AB3A424
= (IA9505001B62C5345479286119EE12C81 [0][41:32] == 10'b01) ? 1'b1 : 1'b0;  generate if (1'b1) begin : I50905559064282CED274D62360FCE175
integer IC12312890F81D79D8CED15EE1E99727F ; always @(posedge ICCFB0F435B37370076102F325BC08D20 or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 )
if (!I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin I6B994CECB5A77B313B1493CB67891E99 <= 1'b0; I109D319C018EB616621364D94266DBCD
<= {64{1'b0}}; IBABAB34D868FD2B2C7A88C42E97BBE11 <= 1'b0; I265478FD9C844733CCACAB4D3F6F7A3F <= 1'b0; IECFDE780B7B9CC7363547C818E204EBB
<= 3'b0; I1B52D4A8BF5D40A682398CBEA678902A <= 11'b0; I9C1F19035765F165886CDE9ADA8857F3 <= 1'b0; I54BE80AB8C90F3E5819921EF5354732A
<= 1'b0; I586C583482F0FD3AF11293684F55AD76 <= 1'b0; I57B81EC60D40AFFA64B92817187C45D7 <= 1'b0; I028038B8A4E4CB73C6DD88AF8C0C9F3E
<= 1'b0; I46B34B7B5B0375E4DD3F84053E6360B7 <= {IE13B4590716ED954FC344B681DC7BBA6 {1'b0}}; I7D0FD152081CEE292550C7730CCA5F75
<= 3'b0; I64D52FE53B2984CB9C38CC7D9230077D <= 11'b0; IE9F53C1FA095EA11A4F2438E8D110DCB <= {IE13B4590716ED954FC344B681DC7BBA6 {1'b0}};
I6EEF1710176D9017BF7C396C5C2DDAD6 <= {IE13B4590716ED954FC344B681DC7BBA6 {1'b0}}; I72AC15FBC2C6EF14364CFFBBB83E3AC0
<= {64{1'b0}}; IFAB2125DC13DFE796F8D4DDBDFC09F4A <= {64{1'b0}}; I9F845E1C893E9E4563815DFDDDFF7E5B <= 1'b0; I674E1FE7EB5BC40955A2009618388E94
<= 1'b0; I2A6B381FD8829A5C8BD04107C91C9378 <= 1'b0; IE68E826F0832B729C0DA0FA2B2697E2E <= 1'b0; I3A905796D2783CA2AD55AEB4DA75441A
<= 1'b0; I1A378769CCB13A524F53158EF54CADD0 <= 1'b0; I5E5A9B8E7ABF32287F37CE45D050FE5F <= 1'b0; I1407533F2D3FCAAA5E6EC4C54A09AEB5
<= 1'b0; IE8B637460BB6B1FB35EB926F2D20C02B <= 1'b0; ID5AB6F130EBFA08B3BFFD3C140B232D7 <= 64'b0; I2D1CB7F5C024D3CED1F017A4D3BC1F55
<= 1'b0; for (IC12312890F81D79D8CED15EE1E99727F = 0; IC12312890F81D79D8CED15EE1E99727F < IE13B4590716ED954FC344B681DC7BBA6 ;
IC12312890F81D79D8CED15EE1E99727F = IC12312890F81D79D8CED15EE1E99727F + 1) IA9505001B62C5345479286119EE12C81 [IC12312890F81D79D8CED15EE1E99727F ]
<= {64{1'b0}}; end else begin I109D319C018EB616621364D94266DBCD <= (I5E5A9B8E7ABF32287F37CE45D050FE5F == 1'b1) ?
I72AC15FBC2C6EF14364CFFBBB83E3AC0 : IFAB2125DC13DFE796F8D4DDBDFC09F4A ; IBABAB34D868FD2B2C7A88C42E97BBE11 <= I9F845E1C893E9E4563815DFDDDFF7E5B
| I2A6B381FD8829A5C8BD04107C91C9378 | I674E1FE7EB5BC40955A2009618388E94 ; I265478FD9C844733CCACAB4D3F6F7A3F <= IE68E826F0832B729C0DA0FA2B2697E2E
| I1A378769CCB13A524F53158EF54CADD0 | I3A905796D2783CA2AD55AEB4DA75441A ; I9C1F19035765F165886CDE9ADA8857F3 <= I5E5A9B8E7ABF32287F37CE45D050FE5F
| I1407533F2D3FCAAA5E6EC4C54A09AEB5 | I3A905796D2783CA2AD55AEB4DA75441A ; I54BE80AB8C90F3E5819921EF5354732A <= I93AE636CE82DE94CB11ACCF59F8C2254 ;
I586C583482F0FD3AF11293684F55AD76 <= (I028038B8A4E4CB73C6DD88AF8C0C9F3E == 1'b1) ? ~IA9505001B62C5345479286119EE12C81 [0][34]
: I586C583482F0FD3AF11293684F55AD76 ; I028038B8A4E4CB73C6DD88AF8C0C9F3E <= I6EEF1710176D9017BF7C396C5C2DDAD6 & I54BE80AB8C90F3E5819921EF5354732A ;
I46B34B7B5B0375E4DD3F84053E6360B7 [0] <= (I6EEF1710176D9017BF7C396C5C2DDAD6 & IE12D7FB0707DA0B72DA8BD64B6FAEFEB
& IDA82F4C78A43B62E1C09ED19A1443221 )| (I46B34B7B5B0375E4DD3F84053E6360B7 [0] & ~IE9F53C1FA095EA11A4F2438E8D110DCB [0]);
IA9505001B62C5345479286119EE12C81 [0] <= I2AED852F071D7FF5A04BEFAF4E7F3B0F ; IE9F53C1FA095EA11A4F2438E8D110DCB [0]
<= I9B9FF20B523F68871F4D27848F9B4E44 ; I6EEF1710176D9017BF7C396C5C2DDAD6 [0] <= I694FF88E6CB22CE905A2A9A9E00AF7F1 ;
I64D52FE53B2984CB9C38CC7D9230077D <= (I028038B8A4E4CB73C6DD88AF8C0C9F3E == 1'b1) ? IA9505001B62C5345479286119EE12C81 [0][50:40]
: I64D52FE53B2984CB9C38CC7D9230077D ; I72AC15FBC2C6EF14364CFFBBB83E3AC0 <= {IA9505001B62C5345479286119EE12C81 [1][7:0],
IA9505001B62C5345479286119EE12C81 [1][15:8], IA9505001B62C5345479286119EE12C81 [1][23:16], IA9505001B62C5345479286119EE12C81 [1][31:24],
IA9505001B62C5345479286119EE12C81 [1][39:32], IA9505001B62C5345479286119EE12C81 [1][47:40], IA9505001B62C5345479286119EE12C81 [1][55:48],
IA9505001B62C5345479286119EE12C81 [1][63:56]}; IFAB2125DC13DFE796F8D4DDBDFC09F4A <= {IA9505001B62C5345479286119EE12C81 [0][39:32],
IA9505001B62C5345479286119EE12C81 [0][47:40], IA9505001B62C5345479286119EE12C81 [0][55:48], IA9505001B62C5345479286119EE12C81 [0][63:56],
IA9505001B62C5345479286119EE12C81 [1][7:0], IA9505001B62C5345479286119EE12C81 [1][15:8], IA9505001B62C5345479286119EE12C81 [1][23:16],
IA9505001B62C5345479286119EE12C81 [1][31:24]}; I9F845E1C893E9E4563815DFDDDFF7E5B <= IE9F53C1FA095EA11A4F2438E8D110DCB [1]
& (I5E5A9B8E7ABF32287F37CE45D050FE5F | (I46B34B7B5B0375E4DD3F84053E6360B7 [1] & ~I5E5A9B8E7ABF32287F37CE45D050FE5F
& ~I586C583482F0FD3AF11293684F55AD76 )); I674E1FE7EB5BC40955A2009618388E94 <= (I7D0FD152081CEE292550C7730CCA5F75
!= 3'b0) ? (IE9F53C1FA095EA11A4F2438E8D110DCB [1] & ~I57B81EC60D40AFFA64B92817187C45D7 ) : 1'b0; I2A6B381FD8829A5C8BD04107C91C9378
<= I049E6CF82F9492802746D564E2B88117 & (I1407533F2D3FCAAA5E6EC4C54A09AEB5 | (I46B34B7B5B0375E4DD3F84053E6360B7 [1]
& ~I1407533F2D3FCAAA5E6EC4C54A09AEB5 & I586C583482F0FD3AF11293684F55AD76 )); IE68E826F0832B729C0DA0FA2B2697E2E <=
I46B34B7B5B0375E4DD3F84053E6360B7 [1] & ~I5E5A9B8E7ABF32287F37CE45D050FE5F & ~I586C583482F0FD3AF11293684F55AD76 ;
I3A905796D2783CA2AD55AEB4DA75441A <= (I7D0FD152081CEE292550C7730CCA5F75 != 3'b0) ? (IE9F53C1FA095EA11A4F2438E8D110DCB [1]
& ~I57B81EC60D40AFFA64B92817187C45D7 ) : 1'b0; I1A378769CCB13A524F53158EF54CADD0 <= I46B34B7B5B0375E4DD3F84053E6360B7 [1]
& ~I1407533F2D3FCAAA5E6EC4C54A09AEB5 & I586C583482F0FD3AF11293684F55AD76 ; I5E5A9B8E7ABF32287F37CE45D050FE5F <=
(I46B34B7B5B0375E4DD3F84053E6360B7 [1] & ~I5E5A9B8E7ABF32287F37CE45D050FE5F & ~I586C583482F0FD3AF11293684F55AD76 )
| (I5E5A9B8E7ABF32287F37CE45D050FE5F & ~I9F845E1C893E9E4563815DFDDDFF7E5B ); I1407533F2D3FCAAA5E6EC4C54A09AEB5 <=
(I46B34B7B5B0375E4DD3F84053E6360B7 [1] & ~I1407533F2D3FCAAA5E6EC4C54A09AEB5 & I586C583482F0FD3AF11293684F55AD76 )
| (I1407533F2D3FCAAA5E6EC4C54A09AEB5 & ~I2A6B381FD8829A5C8BD04107C91C9378 ); IE8B637460BB6B1FB35EB926F2D20C02B <=
(I6EEF1710176D9017BF7C396C5C2DDAD6 [0] & I54BE80AB8C90F3E5819921EF5354732A ) | (IE8B637460BB6B1FB35EB926F2D20C02B
& ~IE9F53C1FA095EA11A4F2438E8D110DCB [1]); for (IC12312890F81D79D8CED15EE1E99727F = 1; IC12312890F81D79D8CED15EE1E99727F
< IE13B4590716ED954FC344B681DC7BBA6 ; IC12312890F81D79D8CED15EE1E99727F = IC12312890F81D79D8CED15EE1E99727F + 1)
begin I46B34B7B5B0375E4DD3F84053E6360B7 [IC12312890F81D79D8CED15EE1E99727F ] <= I46B34B7B5B0375E4DD3F84053E6360B7 [IC12312890F81D79D8CED15EE1E99727F
- 1]; IA9505001B62C5345479286119EE12C81 [IC12312890F81D79D8CED15EE1E99727F ] <= IA9505001B62C5345479286119EE12C81 [IC12312890F81D79D8CED15EE1E99727F
- 1]; IE9F53C1FA095EA11A4F2438E8D110DCB [IC12312890F81D79D8CED15EE1E99727F ] <= IE9F53C1FA095EA11A4F2438E8D110DCB [IC12312890F81D79D8CED15EE1E99727F
- 1]; I6EEF1710176D9017BF7C396C5C2DDAD6 [IC12312890F81D79D8CED15EE1E99727F ] <= I6EEF1710176D9017BF7C396C5C2DDAD6 [IC12312890F81D79D8CED15EE1E99727F
- 1]; end if (I57B81EC60D40AFFA64B92817187C45D7 ) begin if (IE68E826F0832B729C0DA0FA2B2697E2E | I1A378769CCB13A524F53158EF54CADD0
| I3A905796D2783CA2AD55AEB4DA75441A ) begin I6B994CECB5A77B313B1493CB67891E99 <= I586C583482F0FD3AF11293684F55AD76 ;
IECFDE780B7B9CC7363547C818E204EBB <= I7D0FD152081CEE292550C7730CCA5F75 ; I1B52D4A8BF5D40A682398CBEA678902A <= I64D52FE53B2984CB9C38CC7D9230077D ;
end end else begin if (IE9F53C1FA095EA11A4F2438E8D110DCB ) begin IECFDE780B7B9CC7363547C818E204EBB <= I7D0FD152081CEE292550C7730CCA5F75 ;
I1B52D4A8BF5D40A682398CBEA678902A <= I64D52FE53B2984CB9C38CC7D9230077D ; end end if (I6EEF1710176D9017BF7C396C5C2DDAD6
& I54BE80AB8C90F3E5819921EF5354732A ) begin I57B81EC60D40AFFA64B92817187C45D7 <= IDA82F4C78A43B62E1C09ED19A1443221 ;
I028038B8A4E4CB73C6DD88AF8C0C9F3E <= 1'b1; I7D0FD152081CEE292550C7730CCA5F75 <= IA9505001B62C5345479286119EE12C81 [0][15:13];
I2D1CB7F5C024D3CED1F017A4D3BC1F55 <= I0515522FF1EFD23C59D28B8F6AB3A424 ; end if (IE8B637460BB6B1FB35EB926F2D20C02B
| (I6EEF1710176D9017BF7C396C5C2DDAD6 [0] & I54BE80AB8C90F3E5819921EF5354732A )) ID5AB6F130EBFA08B3BFFD3C140B232D7
<= IA9505001B62C5345479286119EE12C81 [0]; end end endgenerate endmodule 
  module IA68D2B0762B11205E05F2AB6538CBB65 #( parameter I0FC86C5872B740D952167BBB632DE33F = 0, parameter IB71844FFA3AB85FEF45EAB4D35395752
= 512, parameter IDB751C3DD512B8355CF27001F983880A = 16, parameter I66C185998F46A7148163982E39BCD296 = "ecp3", parameter
IE33DC83D2AA8913B2CB48378DAF2547A = 32 ) ( input wire ICCFB0F435B37370076102F325BC08D20 , input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 ,
input wire I93AE636CE82DE94CB11ACCF59F8C2254 , input wire [IDB751C3DD512B8355CF27001F983880A - 1:0] I2AED852F071D7FF5A04BEFAF4E7F3B0F ,
input wire I9B9FF20B523F68871F4D27848F9B4E44 , input wire I694FF88E6CB22CE905A2A9A9E00AF7F1 , input wire ID637623B1855D5BBD98CB5D56E107619 ,
output wire IA05976160EBA6DEFAAAA66970A81B32D , output wire [((IDB751C3DD512B8355CF27001F983880A == 16) ? 32 : 64)
- 1:0] IF249B786312150CAA567D0B3F1DC760E , output wire I99A7C01D853D4CD1BF86EA17B055AE82 , output wire IAB7D8322CEA20D7B2FC0EF19A061CB19 ,
output wire I14B85FB28FCEF458E6F9665F2960F9A2 , output wire [$clog2(IB71844FFA3AB85FEF45EAB4D35395752 + 1) - 1:0]
I5F4B958B42F630F4DF0F2B5578E72A4C , output wire [IE33DC83D2AA8913B2CB48378DAF2547A - 1:0] I08C693C25A115282C35BE10561F37009 ,
output wire ID7A2A8B1E9D92B60194D5FAFAAB15208 , output wire IFAF3E1E717F33D0636699473D114FAAC , output wire I89CFFA73C7546481B72B0FB06D799AEE ,
output wire I3E859D8CBD08E747693AC2BA98F2B947 );  localparam integer I36A1B4EB5B5564A6ED7EA4D42856EFB4 = $clog2(IB71844FFA3AB85FEF45EAB4D35395752 );
localparam integer I6B5887A864947F0A024D375AC57C60DE = (IDB751C3DD512B8355CF27001F983880A == 64) ? 66 : 34; localparam
integer I5A3FC4DD94A14DE370E7B95EAB4E36A3 = (IE33DC83D2AA8913B2CB48378DAF2547A == 64) ? 66 : 34; localparam integer
IA4E3C883F66928FBDB89C1DE143D3C01 = (IDB751C3DD512B8355CF27001F983880A == 64) ? 64 : 32; localparam integer I2F8DC10449A1F24468235753BBC3B988
= $clog2((IB71844FFA3AB85FEF45EAB4D35395752 * (IA4E3C883F66928FBDB89C1DE143D3C01 / IE33DC83D2AA8913B2CB48378DAF2547A ))
+ 1);  wire [I6B5887A864947F0A024D375AC57C60DE - 1:0] IC6787F354EA27E7EED18D80DDE370658 ; wire [IE33DC83D2AA8913B2CB48378DAF2547A
- 1:0] I97BAA0787571D1CFEF8C72A952825BA8 ; wire ID07ACEE11131506A08B73834F606CE6C ; wire I03899612613DE8B2DE608F8716710A4E ;
wire I3D497136C8328CC117FE3C0F58AEDBD1 ; wire IB552918C70C5F8374FC906E0C2225F89 ; wire [IA4E3C883F66928FBDB89C1DE143D3C01
- 1:0] IE593D61A89622FBF1D4D61DBF77B0759 ; wire IEB0657AD1CF8431866F1DACFA91DAE9C ; wire I09D474E43198BB26D683E473E35C90C8 ;
wire IA51154D40B341A92D3FF48956FE47EDD ; wire [IA4E3C883F66928FBDB89C1DE143D3C01 - 1:0] I78FE781BC8B5C49E9E0559250B6D4289 ;
wire IA5B0FE243F631FAA054C108CC3F72E10 ; wire I6DF8AFD2D5E8EFB85D4507AC54B8E25C ; wire I7FC89070B58401310300DEAA85090688 ;
wire [I6B5887A864947F0A024D375AC57C60DE - 1:0] I2CA1A324143051A0AFDEFB54659C657C ; wire IE3B28706B7F8094B8D2A6C7E0F5AAB41 ;
wire [I36A1B4EB5B5564A6ED7EA4D42856EFB4 - 1:0] ID6F8558B7CC8FEFCCFC4931DBBD84FBD ; wire [I2F8DC10449A1F24468235753BBC3B988
- 1:0] I47BF20B234CB874608E4590CFA0DBE88 ; wire [I5A3FC4DD94A14DE370E7B95EAB4E36A3 - 1:0] I967C0730B7C51D10FE97AFAB45FC31E4 ;
wire I7DA036F5B0B44A1D5E3EB0237828A810 ; wire [I36A1B4EB5B5564A6ED7EA4D42856EFB4 - 1:0] IC123DE32267CCF513093EB7DB4A4A676 ;
wire I3D3502037CE2D7E5159EAF99BC9BF78D ;  assign IA05976160EBA6DEFAAAA66970A81B32D = IB552918C70C5F8374FC906E0C2225F89 ;
assign IF249B786312150CAA567D0B3F1DC760E = IE593D61A89622FBF1D4D61DBF77B0759 ; assign I99A7C01D853D4CD1BF86EA17B055AE82
= IEB0657AD1CF8431866F1DACFA91DAE9C ; assign IAB7D8322CEA20D7B2FC0EF19A061CB19 = I09D474E43198BB26D683E473E35C90C8 ;
assign I14B85FB28FCEF458E6F9665F2960F9A2 = IA51154D40B341A92D3FF48956FE47EDD ; assign I5F4B958B42F630F4DF0F2B5578E72A4C
= I47BF20B234CB874608E4590CFA0DBE88 ; assign I08C693C25A115282C35BE10561F37009 = I97BAA0787571D1CFEF8C72A952825BA8 ;
assign ID7A2A8B1E9D92B60194D5FAFAAB15208 = ID07ACEE11131506A08B73834F606CE6C ; assign IFAF3E1E717F33D0636699473D114FAAC
= I7DA036F5B0B44A1D5E3EB0237828A810 ; assign I89CFFA73C7546481B72B0FB06D799AEE = I03899612613DE8B2DE608F8716710A4E ;
assign I3E859D8CBD08E747693AC2BA98F2B947 = ~IE3B28706B7F8094B8D2A6C7E0F5AAB41 ;  assign IC6787F354EA27E7EED18D80DDE370658
= {I6DF8AFD2D5E8EFB85D4507AC54B8E25C , IA5B0FE243F631FAA054C108CC3F72E10 , I78FE781BC8B5C49E9E0559250B6D4289 };
assign I3D497136C8328CC117FE3C0F58AEDBD1 = ~I9ED2A9117D3AEAF54CBA7AD69083BCB7 ; assign {I03899612613DE8B2DE608F8716710A4E ,
ID07ACEE11131506A08B73834F606CE6C , I97BAA0787571D1CFEF8C72A952825BA8 } = I967C0730B7C51D10FE97AFAB45FC31E4 ;  generate
if (IA4E3C883F66928FBDB89C1DE143D3C01 == 32) begin : IDF54FF9484E1DFC8C29689596EA8984F assign IB552918C70C5F8374FC906E0C2225F89
= 1'b0; I792C47F7E7D7705A2329EEB04CA92E91 IDD45DEF33DD1E1740F37FA39376216EB ( .ICCFB0F435B37370076102F325BC08D20
(ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .I93AE636CE82DE94CB11ACCF59F8C2254
(I93AE636CE82DE94CB11ACCF59F8C2254 ), .I2AED852F071D7FF5A04BEFAF4E7F3B0F (I2AED852F071D7FF5A04BEFAF4E7F3B0F [15:0]),
.I9B9FF20B523F68871F4D27848F9B4E44 (I9B9FF20B523F68871F4D27848F9B4E44 ), .I694FF88E6CB22CE905A2A9A9E00AF7F1 (I694FF88E6CB22CE905A2A9A9E00AF7F1 ),
.IF249B786312150CAA567D0B3F1DC760E (IE593D61A89622FBF1D4D61DBF77B0759 ), .I99A7C01D853D4CD1BF86EA17B055AE82 (IEB0657AD1CF8431866F1DACFA91DAE9C ),
.IAB7D8322CEA20D7B2FC0EF19A061CB19 (I09D474E43198BB26D683E473E35C90C8 ), .I14B85FB28FCEF458E6F9665F2960F9A2 (IA51154D40B341A92D3FF48956FE47EDD ),
.I528AB843F22B93013A3EAA53871813E4 (I78FE781BC8B5C49E9E0559250B6D4289 ), .I55EF6D8E66D2B56872BA18F8A67DBCC9 (IA5B0FE243F631FAA054C108CC3F72E10 ),
.ICF9485DAA5CD85FD9CF3AB9F6898D8FC (I6DF8AFD2D5E8EFB85D4507AC54B8E25C ), .I3E859D8CBD08E747693AC2BA98F2B947 (I7FC89070B58401310300DEAA85090688 )
); end endgenerate generate if (IA4E3C883F66928FBDB89C1DE143D3C01 == 64) begin : IB567D629A176C50476C16B489433F82B
assign I09D474E43198BB26D683E473E35C90C8 = IA51154D40B341A92D3FF48956FE47EDD ; IB48580D48DC6311D8E12B4626CE243D8
I4C04DB5B9ADB652783A3EE22975D2BB4 ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .I93AE636CE82DE94CB11ACCF59F8C2254 (I93AE636CE82DE94CB11ACCF59F8C2254 ), .I2AED852F071D7FF5A04BEFAF4E7F3B0F
(I2AED852F071D7FF5A04BEFAF4E7F3B0F ), .I9B9FF20B523F68871F4D27848F9B4E44 (I9B9FF20B523F68871F4D27848F9B4E44 ), .I694FF88E6CB22CE905A2A9A9E00AF7F1
(I694FF88E6CB22CE905A2A9A9E00AF7F1 ), .IA05976160EBA6DEFAAAA66970A81B32D (IB552918C70C5F8374FC906E0C2225F89 ), .IF249B786312150CAA567D0B3F1DC760E
(IE593D61A89622FBF1D4D61DBF77B0759 ), .ID7EB8E74BC37FDF7521CAA3A6410AD1C ( ), .I0DE0BA1FE7C719C02C2286C7BB4E82EC
( ), .I22CD4A94B7889ACD9A7D67943BC18F3B ( ), .I4F75D3BA09A515DCAD40830FB24835A7 ( ), .I14B85FB28FCEF458E6F9665F2960F9A2
(IA51154D40B341A92D3FF48956FE47EDD ), .I528AB843F22B93013A3EAA53871813E4 (I78FE781BC8B5C49E9E0559250B6D4289 ), .I55EF6D8E66D2B56872BA18F8A67DBCC9
(IA5B0FE243F631FAA054C108CC3F72E10 ), .ICF9485DAA5CD85FD9CF3AB9F6898D8FC (I6DF8AFD2D5E8EFB85D4507AC54B8E25C ), .I6CE3395345F58F9D860AC549C8AF1473
(I7FC89070B58401310300DEAA85090688 ) ); end endgenerate pmi_ram_dp # ( .pmi_wr_addr_depth (IB71844FFA3AB85FEF45EAB4D35395752 ),
.pmi_wr_addr_width (I36A1B4EB5B5564A6ED7EA4D42856EFB4 ), .pmi_wr_data_width (I6B5887A864947F0A024D375AC57C60DE ),
.pmi_rd_addr_depth (IB71844FFA3AB85FEF45EAB4D35395752 ), .pmi_rd_addr_width (I36A1B4EB5B5564A6ED7EA4D42856EFB4 ),
.pmi_rd_data_width (I6B5887A864947F0A024D375AC57C60DE ), .pmi_regmode ("reg"), .pmi_family (I66C185998F46A7148163982E39BCD296 ),
.module_type ("pmi_ram_dp") ) I25719AD8557B4584865155DAE07C7840 ( .Data (IC6787F354EA27E7EED18D80DDE370658 ), .RdAddress
(ID6F8558B7CC8FEFCCFC4931DBBD84FBD ), .RdClockEn (1'b1), .RdClock (ICCFB0F435B37370076102F325BC08D20 ), .Reset (I3D497136C8328CC117FE3C0F58AEDBD1 ),
.WE (I3D3502037CE2D7E5159EAF99BC9BF78D ), .WrAddress (IC123DE32267CCF513093EB7DB4A4A676 ), .WrClockEn (1'b1), .WrClock
(ICCFB0F435B37370076102F325BC08D20 ), .Q (I2CA1A324143051A0AFDEFB54659C657C ) ); I6B46C5BDF6C2841AE2EEF22D18B3C8B9
# ( .I61D0345D311EC6FFC08DDDECE5F6127A (IB71844FFA3AB85FEF45EAB4D35395752 ), .I5C6C6CD7723900C21B3A76E887CEE164
(IA4E3C883F66928FBDB89C1DE143D3C01 ), .I64BB723AC8F87F7AEBA73BF190ED5F8F (IE33DC83D2AA8913B2CB48378DAF2547A ), .I846B877ED5AEDADF389E2082E674F6A2
(2) ) I5B7A19877C7417CDB4387DF988625F8B ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ),
.I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .I1A61D2CA45ECC28270C28826CD87FEC3 (I2CA1A324143051A0AFDEFB54659C657C ),
.IC79EC9A9F373F4B71374BDF6EDD31DE6 (1'b0), .I3DAC0A14B4001DD3A76D99313964C3AA (1'b0), .IFF897FEF3F69926A750D8217ADD6AE1C
(ID637623B1855D5BBD98CB5D56E107619 ), .I22B24791BA0E7AA2C686B1B2D776C636 (I7FC89070B58401310300DEAA85090688 ), .I79D313D86841E5141E7629EA606D7AE9
(ID6F8558B7CC8FEFCCFC4931DBBD84FBD ), .I11CEFC90537A67CD1FF01400245362F2 (), .ID7FCE45A65ADDB17F91F73A1B506BB5B
(I47BF20B234CB874608E4590CFA0DBE88 ), .I125028C7446331521D0434C10E8B0007 (I967C0730B7C51D10FE97AFAB45FC31E4 ), .I8BB939FF2AFDE7B2A1E480DCB61CE354
(IE3B28706B7F8094B8D2A6C7E0F5AAB41 ), .I41C63F948E534C7ED9F2471A44C922B2 (), .I07E2A2E89C25B45C36871FC0931EC8EF
(I7DA036F5B0B44A1D5E3EB0237828A810 ), .I38B1AC532E13E69B05492C67EC7070BB (IC123DE32267CCF513093EB7DB4A4A676 ), .I705C64753A50CDA034B5ACB332D71768
(), .I102322A55721851004CB8E1F6AB50BDE (I3D3502037CE2D7E5159EAF99BC9BF78D ), .I233E0C0C8E5150F0CD8258F276D93942
(), .IBE0D6810EBD63B5C428623C578CF6D3A (), .I115E90220158F08B0465E99D7F2561D3 () ); endmodule 
  module I4CACC63B64035D749DE3C4BCF79F626C #( parameter IA0709F456132ABB4EB324E1598AAB825 = 512, parameter IFC796EA7F9507A2288E499F7B9ECC63E
= 512, parameter IDB9D60794264C5F8E5363941194A797B = 3, parameter I50AC25E9687F891BB7188EED025C1323 = 0, parameter
ID7C7F9F2E39BEBEE2ACFA8040034E48D = 16 ) ( input wire ICCFB0F435B37370076102F325BC08D20 , input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 ,
input wire I69B8FD7561F9CA8AAF4E50C5B2DCF850 , input wire IA85D446CD214F6B3CE6418205432D870 , input wire IBB8FE5B389C0BD7BA64F2E05FCDC4485 ,
input wire I45A8F29589769D54C9D702481065CB45 , input wire [7:0] IFF5E23C5A17BB678C108274E28C56424 , input wire [4:0]
IDE425A12275C43D9056DCF647A2D8258 , input wire [2:0] I65B14714ECFCC218D3A788DF7696216B , input wire [2:0] IA1F0CBEC8E9EAD83D0098DD96A1EFC32 ,
input wire IFC18758E8987A9913FD94A5DFEE774E2 , input wire IF5E7E4E58741BF3FE58442AB377ED57F , input wire IF5B4924BEAEA6935367AC2739021882F ,
input wire I7985A5A43CBBBC8E0D3FCFEE38DDF221 , input wire [IDB9D60794264C5F8E5363941194A797B - 1:0] I7E600D684E83043922C1FE27CC6213E4 ,
input wire I93AE636CE82DE94CB11ACCF59F8C2254 , input wire [7:0] I9119CE851F731CBC5834D0370CCA6908 , input wire [$clog2(IA0709F456132ABB4EB324E1598AAB825
+ 1) - 1:0] I9F3623AEB414A15CECD2A8FD8791C79D , input wire [31:0] I36824F33FF142FDE2AFE9BC4759DB690 , input wire
I5E84ED10AD623502BC750C5E797D1428 , input wire IA886199C0F7609B072DAE171DFC98CD8 , input wire IA067043029572C8598E352E0A66EA337 ,
input wire [$clog2(IFC796EA7F9507A2288E499F7B9ECC63E + 1) - 1:0] ICB518A59CAE27DDB6398AB22F5D74259 , input wire
I9F4F7E2C4A4A8FB2780021EDF6E4ADEF , input wire I07B0EBE8FBC21BDBE894D73C90EDC5AB , input wire I44B3CB0FFE4214C92C98CD6ECFC52D5A ,
input wire [31:0] I3D6C771D05CA1A769E61302C086494B8 , output wire [7:0] IC2E260CA356C994048CCB108C7E359D1 , output
wire [7:0] IE707B5D4A74BA1BD745B52E0C07932C0 , output wire I6E70C748D9C56227AB1182F36658AE5C , output wire I59B23598E8ADE1982F184EF67BEB0979 ,
output wire I33E409903692F5ECA2EC3553F9D1659E , output wire I437E57D42FB91B674CCBCC915BF9D653 , output wire I55AFDDE17B53D7F65849D39B02B07417 ,
output wire [31:0] I65FE2DB4E1CB5A488A45D60041AB5F64 , output wire [63:0] I0C796C206FE7060B578156D0110461EB , output
wire IFC86A6522A8CA080A0DB7F384D9CE6FA , output wire I484F77D7967D25736EB27A0ED76CCB5F , output wire I7E0431D7F1A92C0ED1F030F36BF809B7 ,
output wire I3E6965EC606FD6C2871F2C0993204C57 , output wire IFF25B820DFD457D71B32B130ABE5DA3F , output wire I20FA57C9A87CB2AA26088D9FA1743F70 ,
output wire I51C881E8B9B36D7A724BC7B8EC533957 , output wire [7:0] ID3E7F4B58943229FEE6313A36B3F8693 , output wire
[4:0] I1FDEC1735547330C00A0B8DFE1FB10C3 , output wire [2:0] IBD6A65D48B4A68CA0D2A82F79053757B , output wire I15EC78E3DE1101BFF2B227962683E113 ,
output wire [31:0] I7C4DADE2C05F6DCECCAF7AD6F7BF2FF8 , output wire IEEFA85D6664F09687B5CA591C701DC34 , output wire
ID4A284C76C6EABEEBA8E0AE18003FBAC , output wire I6010C20131B976554A498745FEEEB580 , output wire [ID7C7F9F2E39BEBEE2ACFA8040034E48D
- 1:0] I46E8CA15DC1E8B3B2200999A53029704 , output wire [1:0] IEC45B60C7D1A49FFA84D3F5D121A2579 , output wire [2:0]
I9AF46E2AA924FA7E0F5D7290324BABF9 , output wire I59D9A9A677978229C1F87AA1A3A0C304 , output wire I9301CE4E9B877D08EDBD1584D6BE017A ,
output wire I51698892CBD372EE66AF3EA4D0ECE23F , output wire I1347408C9E757F34EA4D78F53447BD9B , output wire [IDB9D60794264C5F8E5363941194A797B
- 1:0] I2BE88607F3C31B47400F3A35E08B7EAD , output wire [31:0] I7D901091F9E0741061C75B54467D48A0 , output wire I7AEBDB3D2CD4891A528BA81F5F54B20D ,
output wire [10:0] ID16819FEAA95700005E383E7DA0C8E13 , output wire [3:0] IE0337CA803FBA20F38A0CD2A900C6534 , output
wire [3:0] I592A6A3BA99B09C24695C7A609F9053F , output wire [3:0] I40EF39BB4F4F4A031C8FD1026EF53063 , output wire
I42427E866FF31BC28E35C71EC172E26B , output wire I368749E68EAF9F462385FAD36180A9FE ); `include "pcisig_constants.v"
`include "wishbone_utils.v"
 localparam I15DA3B10E1E0658D2D01B744DF560903 = 3; localparam I1797388B2E6E3CB5EE600DD85605F982 = $clog2(I15DA3B10E1E0658D2D01B744DF560903 );
localparam IDE267FF256F75C9698907411CE334A5B = $clog2(IA0709F456132ABB4EB324E1598AAB825 + 1); localparam I30AF2C9FF2EEDF02869CDAC1AAC433BC
= $clog2(IFC796EA7F9507A2288E499F7B9ECC63E + 1); localparam I3662C12143A4A1B904AC8798CEEF0125 = 5'b00000, I257DF24B77C5CA85F676E7FFA065CE94
= 5'b00001, I54DD54FD7FB944705CE08C2B291B87A7 = 5'b00010, I962A83F6AB78F0114DD9D85409B29E8F = 5'b00011, IA4997CC969740D4CF1FC8E4E9C2B5DA7
= 5'b00100, I8EBFD17705709FF6F2CAA85EA87D66D4 = 5'b00101, I56AC73D28E70D2F78200164359CC0E9A = 5'b00110, I499DB4E92AEE1C97FE024F6FD8CDEB8A
= 5'b00111, IABEE3580E02F366EC5560A9CFC5CC953 = 5'b01000, I2D358EAE916810B434B6C76F7C7C5673 = 5'b01001, I174E152AA0198C30C57B401C947D37C1
= 5'b01010, I3C15F904BACDB851EFC4C548820E98B8 = 5'b01011, I61A7D75570E89738696B9598A883C1CD = 5'b01100, I29C10DD8DAC8AB31273614BA27A5E29C
= 5'b01101, IF5A7A7CE92502E2DF9F0601605A38637 = 5'b01110, I5021A214EB457E909E76C621F6DD12B1 = 5'b01111, IFAC7B411ECB5421590DDAA0B7B34F238
= 5'b10000, I248DCDE6260EE21AB43E9E1EF6D603EF = 5'b10001, IC495D10CCC7452A18D769BDD99794652 = 5'b10010, IEAE55E29AC7D8EC5093BF4C91D5CFFCE
= 5'b10011, I6EA1237B063AFA6C82E354D0001BEF41 = 5'b10100, ID1D4A1F29119D84947D94DCCD5BDF6A9 = 5'b10101, IF86E23BE5E6D56399363666A2BDC7A6A
= 5'b10110, I264B836E51E7F23F603A59DFDC8D2C8A = 5'b10111, I05E305FFF5B6CDE122F8935EE521D523 = 5'b11000, IFE8FF815A0D8FDD4B9426B3849E23E02
= 5'b11001;  reg [3:0] I11FD35FED78BCB8861FACB9A1E3A4C35 ; reg [3:0] IC52F3B77F7E45A74323561D6A6F6028A ; reg I0FF03F7D70F3047C91A55F9744DDD7AE ;
reg [11:0] IAC85A6B0EE1F3079B60C115CB476DF06 ; reg [8:0] I71DBDE411F9CED520FD43A4EF5CBD656 ; reg [7:0] IBFF7FD594C616C9EBAD12448149DA576 ;
reg I0C9CC98CD774EDC9DF9AB513E5A8FB57 ; reg I26F46DF735C89C3DA76F7F404A5F650F ; reg [7:0] I5AF6C20F3950D58007B9C0BEA7C87198 ;
reg I533559C7D3A6FC7D4A2E49A02AFC9137 ; reg IF9A51F60DF053D68A5D57FECB5AB7ACB ; reg I916551CA30E7A94681BA2B3415BF85FA ;
reg I4A3B5CD6A0CBD18332DCF8ECB309CC92 ; reg [31:0] I2931854F66F4E6D5E96ED7D73266F38E ; reg [I1797388B2E6E3CB5EE600DD85605F982
- 1:0] IDA48F17DCE4BB1F6A04CBB23CCB4C3A5 ; reg IC93C4C87277AF77C73E35A77E14FC4B1 ; reg I54BE80AB8C90F3E5819921EF5354732A ;
reg I623116EB4A13517E3733A1778B496560 ; reg I511F58CE0ACA83EE959D1BF6C4EAFA7F ; reg [7:0] I7E9516402D6933186513EB5B37336278 ;
reg [4:0] IA1EA4D4C05E159614ABC1E6D9CABE3BB ; reg [2:0] I8916D921407646CE03BABA39B922EE09 ; reg I7FA4C54BD6B551C794EE0EA588CBD4C7 ;
reg I9C46AA186B65717669AB8B1F7ED02022 ; reg IE4E0DDAB16DD8E970672626428251866 ; reg IE12D7FB0707DA0B72DA8BD64B6FAEFEB ;
reg I15C3BE43949B828A0A578329FE2EDE6B ; reg IE655D625D2EB067AC17967E600BE5FBD ; reg IABBE7E409672B3D3CE209351AE63C530 ;
reg I9962CDA8EE94C7BDFB23FE70815056E4 ; reg I7732946249B5963DFD9C95EC611A1D2C ; reg [6:0] I54D7451A32675B2129629BC41778D6D6 ;
reg [4:0] I8AC99AB880823B01C00D137F89AABEF8 ; reg [4:0] IF15E5692F18C2355720A228228564D0B ; reg I9B8138DCE156F7C31EB5914EF01F183C ;
reg [7:0] IB9A23596C80981B9B1CF7E12A76E71AC ; reg [4:0] I288715DFB3893A064D51571152559F12 ; reg [2:0] I86B9557FA0123B8105E34300F4FCD447 ;
reg [IDE267FF256F75C9698907411CE334A5B - 1:0] I3EC90F87E70407C2A46DA25A8CA9065B ; reg [31:0] I9E40C3A9F9E3CDFC05F95566701DFB02 ;
reg ICFC6D424C8D5969FAC575FE0538F20F3 ; reg ICDFF33095CB0890DA2F167B63251EC67 ; reg IEDEC097EECBEE6B592219F6FEFFC7C2A ;
reg [10:0] I9E185DF5B08D79D1F56FD64627570AE0 ; reg I08AAFC572BC9A693B4E7C04DFD77FEAF ; reg [7:0] I0C9005A5E5456704CE9C506A03373402 ;
reg [IDB9D60794264C5F8E5363941194A797B - 1:0] I5B0AA124C4ADA63A064AF2CAFA1098FD ; reg [3:0] I93F6D99D18FD6FF40EF5AD5288D5C88E ;
reg [63:0] I83F18730E4735495B20E29C862E672F1 ; reg [13:0] I18D210808E8E4FD4E19269D50B767EF6 ; reg [10:0] I84B10D95B4B5E01F827E0D4D81BF476B ;
reg [7:0] I539C1D01FC349447001EB93E17D37611 ; reg [31:0] I2C5E6805594DFF3B9EB915045ABF7575 ; reg [I30AF2C9FF2EEDF02869CDAC1AAC433BC
- 1:0] I909A2BB1C99AC88EE130F2C2B36CD5AB ; reg I893DF0D582AF0617B44879E65C202360 ; reg I2967174B668E2BB5A635A3F85DFF312B ;
reg I2212D954BC70C49C1F608E169DC873BC ; reg I5B3BB6CF473F793585E2668A9A7136C8 ; reg [ID7C7F9F2E39BEBEE2ACFA8040034E48D
- 1:0] IC7779D4175ADF3F75C21392F9E824B6D ; reg [1:0] IA6B00370F90E5BFE7B5D8852390CF107 ; reg [2:0] I369C3845EEBC3367BADAF446789A185D ;
reg I57E5F0C022683CA716D05ABE3408A469 ; reg IE7D8E2A0B7B7689804FFDF702BF724A6 ; reg I6F3C14B2AF4F4232F642DBEB36DCF09E ;
reg I33F9C80AA280FFCBE2A2CB54C2056CC5 ; reg [IDB9D60794264C5F8E5363941194A797B - 1:0] I5A4554E3FF0F3BAFC519CDF46237B987 ;
reg [31:0] I074FD9C5AE408613B3750B75A6125486 ; reg I0EBD58BCF1D55F648B20B722C25EA4A8 ; reg [10:0] I30D7DB78C2B62A00872F044F1A2F39A2 ;
reg [10:0] IA934CBE3CC9AEBA0C32AA4C7EFA4954C ; reg [3:0] I13C229A5BDE90D9F920D8F4D218106DE ; reg I037773E6A298229B4A19627ABA272E81 ;
reg I36FECBB048E15937DC767259CBABEDCB ; wire [7:0] IC4C940842A3072C3A9C40616C6A213F2 ; wire [4:0] IE8010EDEC4159FBD688A550900D0006D ;
wire [2:0] I6345C4C803C15670FB2665AEA7AA4E33 ; wire IDEA2A0E5DD71C950358A21DDB6565B0A ; wire I93FEA934E2F91A4D5E773376B9B26FED ;
wire [31:0] I44109A75F9883AA09218902DA5B2CBB3 ;  assign IC2E260CA356C994048CCB108C7E359D1 = IBFF7FD594C616C9EBAD12448149DA576 ;
assign IE707B5D4A74BA1BD745B52E0C07932C0 = I5AF6C20F3950D58007B9C0BEA7C87198 ; assign I6E70C748D9C56227AB1182F36658AE5C
= I0C9CC98CD774EDC9DF9AB513E5A8FB57 ; assign I59B23598E8ADE1982F184EF67BEB0979 = I26F46DF735C89C3DA76F7F404A5F650F ;
assign I33E409903692F5ECA2EC3553F9D1659E = I533559C7D3A6FC7D4A2E49A02AFC9137 ; assign I437E57D42FB91B674CCBCC915BF9D653
= IF9A51F60DF053D68A5D57FECB5AB7ACB ; assign I55AFDDE17B53D7F65849D39B02B07417 = I4A3B5CD6A0CBD18332DCF8ECB309CC92 ;
assign I65FE2DB4E1CB5A488A45D60041AB5F64 = {I2931854F66F4E6D5E96ED7D73266F38E [7:0], I2931854F66F4E6D5E96ED7D73266F38E [15:8],
I2931854F66F4E6D5E96ED7D73266F38E [23:16], I2931854F66F4E6D5E96ED7D73266F38E [31:24]}; assign I0C796C206FE7060B578156D0110461EB
= I83F18730E4735495B20E29C862E672F1 ; assign IFC86A6522A8CA080A0DB7F384D9CE6FA = IE12D7FB0707DA0B72DA8BD64B6FAEFEB ;
assign I484F77D7967D25736EB27A0ED76CCB5F = I9C46AA186B65717669AB8B1F7ED02022 ; assign I7E0431D7F1A92C0ED1F030F36BF809B7
= IE4E0DDAB16DD8E970672626428251866 ; assign I3E6965EC606FD6C2871F2C0993204C57 = I15C3BE43949B828A0A578329FE2EDE6B ;
assign IFF25B820DFD457D71B32B130ABE5DA3F = IE655D625D2EB067AC17967E600BE5FBD ; assign I20FA57C9A87CB2AA26088D9FA1743F70
= IABBE7E409672B3D3CE209351AE63C530 ; assign I51C881E8B9B36D7A724BC7B8EC533957 = I511F58CE0ACA83EE959D1BF6C4EAFA7F ;
assign ID3E7F4B58943229FEE6313A36B3F8693 = I7E9516402D6933186513EB5B37336278 ; assign I1FDEC1735547330C00A0B8DFE1FB10C3
= IA1EA4D4C05E159614ABC1E6D9CABE3BB ; assign IBD6A65D48B4A68CA0D2A82F79053757B = I8916D921407646CE03BABA39B922EE09 ;
assign I15EC78E3DE1101BFF2B227962683E113 = IEDEC097EECBEE6B592219F6FEFFC7C2A ; assign I7C4DADE2C05F6DCECCAF7AD6F7BF2FF8
= I2C5E6805594DFF3B9EB915045ABF7575 ; assign IEEFA85D6664F09687B5CA591C701DC34 = I893DF0D582AF0617B44879E65C202360 ;
assign ID4A284C76C6EABEEBA8E0AE18003FBAC = I2212D954BC70C49C1F608E169DC873BC ; assign I6010C20131B976554A498745FEEEB580
= I5B3BB6CF473F793585E2668A9A7136C8 ; assign I46E8CA15DC1E8B3B2200999A53029704 = IC7779D4175ADF3F75C21392F9E824B6D ;
assign IEC45B60C7D1A49FFA84D3F5D121A2579 = IA6B00370F90E5BFE7B5D8852390CF107 ; assign I9AF46E2AA924FA7E0F5D7290324BABF9
= I369C3845EEBC3367BADAF446789A185D ; assign I59D9A9A677978229C1F87AA1A3A0C304 = I57E5F0C022683CA716D05ABE3408A469 ;
assign I9301CE4E9B877D08EDBD1584D6BE017A = IE7D8E2A0B7B7689804FFDF702BF724A6 ; assign I51698892CBD372EE66AF3EA4D0ECE23F
= I6F3C14B2AF4F4232F642DBEB36DCF09E ; assign I1347408C9E757F34EA4D78F53447BD9B = I33F9C80AA280FFCBE2A2CB54C2056CC5 ;
assign I2BE88607F3C31B47400F3A35E08B7EAD = I5A4554E3FF0F3BAFC519CDF46237B987 ; assign I7D901091F9E0741061C75B54467D48A0
= {I074FD9C5AE408613B3750B75A6125486 [7:0], I074FD9C5AE408613B3750B75A6125486 [15:8], I074FD9C5AE408613B3750B75A6125486 [23:16],
I074FD9C5AE408613B3750B75A6125486 [31:24]}; assign I7AEBDB3D2CD4891A528BA81F5F54B20D = I0EBD58BCF1D55F648B20B722C25EA4A8 ;
assign ID16819FEAA95700005E383E7DA0C8E13 = I30D7DB78C2B62A00872F044F1A2F39A2 ; assign IE0337CA803FBA20F38A0CD2A900C6534
= I11FD35FED78BCB8861FACB9A1E3A4C35 ; assign I592A6A3BA99B09C24695C7A609F9053F = IC52F3B77F7E45A74323561D6A6F6028A ;
assign I40EF39BB4F4F4A031C8FD1026EF53063 = I13C229A5BDE90D9F920D8F4D218106DE ; assign I42427E866FF31BC28E35C71EC172E26B
= I037773E6A298229B4A19627ABA272E81 ; assign I368749E68EAF9F462385FAD36180A9FE = I36FECBB048E15937DC767259CBABEDCB ;
 assign IC4C940842A3072C3A9C40616C6A213F2 = (I511F58CE0ACA83EE959D1BF6C4EAFA7F & I9C46AA186B65717669AB8B1F7ED02022 )
? I7E9516402D6933186513EB5B37336278 : IFF5E23C5A17BB678C108274E28C56424 ; assign IE8010EDEC4159FBD688A550900D0006D
= (I511F58CE0ACA83EE959D1BF6C4EAFA7F & I9C46AA186B65717669AB8B1F7ED02022 ) ? IA1EA4D4C05E159614ABC1E6D9CABE3BB :
IDE425A12275C43D9056DCF647A2D8258 ; assign I6345C4C803C15670FB2665AEA7AA4E33 = (I511F58CE0ACA83EE959D1BF6C4EAFA7F
& I9C46AA186B65717669AB8B1F7ED02022 ) ? I8916D921407646CE03BABA39B922EE09 : I65B14714ECFCC218D3A788DF7696216B ;
assign IDEA2A0E5DD71C950358A21DDB6565B0A = (I7E600D684E83043922C1FE27CC6213E4 ) ? 1'b1 : 1'b0; assign I93FEA934E2F91A4D5E773376B9B26FED
= (I9C46AA186B65717669AB8B1F7ED02022 & IF5E7E4E58741BF3FE58442AB377ED57F ) | (IE12D7FB0707DA0B72DA8BD64B6FAEFEB
& IFC18758E8987A9913FD94A5DFEE774E2 ) | (IE4E0DDAB16DD8E970672626428251866 & IF5B4924BEAEA6935367AC2739021882F )
| ((I15C3BE43949B828A0A578329FE2EDE6B | IE655D625D2EB067AC17967E600BE5FBD ) & IDEA2A0E5DD71C950358A21DDB6565B0A )
| (IABBE7E409672B3D3CE209351AE63C530 & I7985A5A43CBBBC8E0D3FCFEE38DDF221 ); assign I44109A75F9883AA09218902DA5B2CBB3
= {I3D6C771D05CA1A769E61302C086494B8 [7:0], I3D6C771D05CA1A769E61302C086494B8 [15:8], I3D6C771D05CA1A769E61302C086494B8 [23:16],
I3D6C771D05CA1A769E61302C086494B8 [31:24]};  always @(*) begin IF15E5692F18C2355720A228228564D0B = I8AC99AB880823B01C00D137F89AABEF8 ;
case (I8AC99AB880823B01C00D137F89AABEF8 ) I3662C12143A4A1B904AC8798CEEF0125 : begin if (I9F3623AEB414A15CECD2A8FD8791C79D
> 2) IF15E5692F18C2355720A228228564D0B = I257DF24B77C5CA85F676E7FFA065CE94 ; end I257DF24B77C5CA85F676E7FFA065CE94
: begin if (IA886199C0F7609B072DAE171DFC98CD8 == 1'b1) IF15E5692F18C2355720A228228564D0B = I54DD54FD7FB944705CE08C2B291B87A7 ;
end I54DD54FD7FB944705CE08C2B291B87A7 : begin IF15E5692F18C2355720A228228564D0B = I962A83F6AB78F0114DD9D85409B29E8F ;
end I962A83F6AB78F0114DD9D85409B29E8F : begin IF15E5692F18C2355720A228228564D0B = IA4997CC969740D4CF1FC8E4E9C2B5DA7 ;
end IA4997CC969740D4CF1FC8E4E9C2B5DA7 : begin if (I623116EB4A13517E3733A1778B496560 ) IF15E5692F18C2355720A228228564D0B
= I56AC73D28E70D2F78200164359CC0E9A ; else IF15E5692F18C2355720A228228564D0B = I8EBFD17705709FF6F2CAA85EA87D66D4 ;
end I8EBFD17705709FF6F2CAA85EA87D66D4 : begin if (ICFC6D424C8D5969FAC575FE0538F20F3 ) IF15E5692F18C2355720A228228564D0B
= I56AC73D28E70D2F78200164359CC0E9A ; end I56AC73D28E70D2F78200164359CC0E9A : begin if (IDA48F17DCE4BB1F6A04CBB23CCB4C3A5
== 0) IF15E5692F18C2355720A228228564D0B = I499DB4E92AEE1C97FE024F6FD8CDEB8A ; end I499DB4E92AEE1C97FE024F6FD8CDEB8A
: begin if (I93FEA934E2F91A4D5E773376B9B26FED ) if (I9962CDA8EE94C7BDFB23FE70815056E4 ) IF15E5692F18C2355720A228228564D0B
= IC495D10CCC7452A18D769BDD99794652 ; else if (I511F58CE0ACA83EE959D1BF6C4EAFA7F ) IF15E5692F18C2355720A228228564D0B
= IABEE3580E02F366EC5560A9CFC5CC953 ; else IF15E5692F18C2355720A228228564D0B = I2D358EAE916810B434B6C76F7C7C5673 ;
else IF15E5692F18C2355720A228228564D0B = IFAC7B411ECB5421590DDAA0B7B34F238 ; end IABEE3580E02F366EC5560A9CFC5CC953
: begin if (ICDFF33095CB0890DA2F167B63251EC67 ) IF15E5692F18C2355720A228228564D0B = I2D358EAE916810B434B6C76F7C7C5673 ;
end I2D358EAE916810B434B6C76F7C7C5673 : begin  IF15E5692F18C2355720A228228564D0B = I174E152AA0198C30C57B401C947D37C1 ;
end I174E152AA0198C30C57B401C947D37C1 : begin if (I511F58CE0ACA83EE959D1BF6C4EAFA7F ) begin if (IA886199C0F7609B072DAE171DFC98CD8
== 1'b1) IF15E5692F18C2355720A228228564D0B = I29C10DD8DAC8AB31273614BA27A5E29C ; end else IF15E5692F18C2355720A228228564D0B
= I3C15F904BACDB851EFC4C548820E98B8 ; end I3C15F904BACDB851EFC4C548820E98B8 : begin if (I07B0EBE8FBC21BDBE894D73C90EDC5AB
& (IA934CBE3CC9AEBA0C32AA4C7EFA4954C == 1)) IF15E5692F18C2355720A228228564D0B = IF5A7A7CE92502E2DF9F0601605A38637 ;
end I29C10DD8DAC8AB31273614BA27A5E29C : begin if (I07B0EBE8FBC21BDBE894D73C90EDC5AB & (IA934CBE3CC9AEBA0C32AA4C7EFA4954C
== 1)) IF15E5692F18C2355720A228228564D0B = IF5A7A7CE92502E2DF9F0601605A38637 ; end IF5A7A7CE92502E2DF9F0601605A38637
: begin IF15E5692F18C2355720A228228564D0B = I5021A214EB457E909E76C621F6DD12B1 ; end I5021A214EB457E909E76C621F6DD12B1
: begin if (I7FA4C54BD6B551C794EE0EA588CBD4C7 ) IF15E5692F18C2355720A228228564D0B = I05E305FFF5B6CDE122F8935EE521D523 ;
else if (I50AC25E9687F891BB7188EED025C1323 ) IF15E5692F18C2355720A228228564D0B = IFE8FF815A0D8FDD4B9426B3849E23E02 ;
else IF15E5692F18C2355720A228228564D0B = I3662C12143A4A1B904AC8798CEEF0125 ; end I05E305FFF5B6CDE122F8935EE521D523
: begin if (I9F4F7E2C4A4A8FB2780021EDF6E4ADEF ) if (I50AC25E9687F891BB7188EED025C1323 ) IF15E5692F18C2355720A228228564D0B
= IFE8FF815A0D8FDD4B9426B3849E23E02 ; else IF15E5692F18C2355720A228228564D0B = I3662C12143A4A1B904AC8798CEEF0125 ;
end IFAC7B411ECB5421590DDAA0B7B34F238 : begin if (I511F58CE0ACA83EE959D1BF6C4EAFA7F ) begin if (ICDFF33095CB0890DA2F167B63251EC67 )
IF15E5692F18C2355720A228228564D0B = I248DCDE6260EE21AB43E9E1EF6D603EF ; end else begin if (I9962CDA8EE94C7BDFB23FE70815056E4 )
IF15E5692F18C2355720A228228564D0B = I6EA1237B063AFA6C82E354D0001BEF41 ; else IF15E5692F18C2355720A228228564D0B =
IF5A7A7CE92502E2DF9F0601605A38637 ; end end I248DCDE6260EE21AB43E9E1EF6D603EF : begin if (I08AAFC572BC9A693B4E7C04DFD77FEAF
== 1'b1) if (I9962CDA8EE94C7BDFB23FE70815056E4 )  IF15E5692F18C2355720A228228564D0B = I6EA1237B063AFA6C82E354D0001BEF41 ;
else IF15E5692F18C2355720A228228564D0B = IF5A7A7CE92502E2DF9F0601605A38637 ; end IC495D10CCC7452A18D769BDD99794652
: begin if (ICB518A59CAE27DDB6398AB22F5D74259 > 2) IF15E5692F18C2355720A228228564D0B = I6EA1237B063AFA6C82E354D0001BEF41 ;
end IEAE55E29AC7D8EC5093BF4C91D5CFFCE : begin if (I2967174B668E2BB5A635A3F85DFF312B ) IF15E5692F18C2355720A228228564D0B
= I2D358EAE916810B434B6C76F7C7C5673 ; end I6EA1237B063AFA6C82E354D0001BEF41 : begin IF15E5692F18C2355720A228228564D0B
= ID1D4A1F29119D84947D94DCCD5BDF6A9 ; end ID1D4A1F29119D84947D94DCCD5BDF6A9 : begin IF15E5692F18C2355720A228228564D0B
= IF86E23BE5E6D56399363666A2BDC7A6A ; end IF86E23BE5E6D56399363666A2BDC7A6A : begin IF15E5692F18C2355720A228228564D0B
= I264B836E51E7F23F603A59DFDC8D2C8A ; end I264B836E51E7F23F603A59DFDC8D2C8A : begin if (I7732946249B5963DFD9C95EC611A1D2C )
IF15E5692F18C2355720A228228564D0B = IF5A7A7CE92502E2DF9F0601605A38637 ; else if (I511F58CE0ACA83EE959D1BF6C4EAFA7F )
IF15E5692F18C2355720A228228564D0B = IABEE3580E02F366EC5560A9CFC5CC953 ; else IF15E5692F18C2355720A228228564D0B =
IEAE55E29AC7D8EC5093BF4C91D5CFFCE ; end IFE8FF815A0D8FDD4B9426B3849E23E02 : begin if (~IEDEC097EECBEE6B592219F6FEFFC7C2A
& ~(|I0C9005A5E5456704CE9C506A03373402 )) IF15E5692F18C2355720A228228564D0B = I3662C12143A4A1B904AC8798CEEF0125 ;
end default : begin end endcase end  always @(posedge ICCFB0F435B37370076102F325BC08D20 or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 )
begin : I50905559064282CED274D62360FCE175 if (~I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin I11FD35FED78BCB8861FACB9A1E3A4C35
<= 4'hf; IC52F3B77F7E45A74323561D6A6F6028A <= 4'hf; I0FF03F7D70F3047C91A55F9744DDD7AE <= 1'b0; IAC85A6B0EE1F3079B60C115CB476DF06
<= 12'b0; I71DBDE411F9CED520FD43A4EF5CBD656 <= 9'b0; IBFF7FD594C616C9EBAD12448149DA576 <= 8'b0; I0C9CC98CD774EDC9DF9AB513E5A8FB57
<= 1'b0; I26F46DF735C89C3DA76F7F404A5F650F <= 1'b0; I5AF6C20F3950D58007B9C0BEA7C87198 <= 8'b0; I533559C7D3A6FC7D4A2E49A02AFC9137
<= 1'b0; IF9A51F60DF053D68A5D57FECB5AB7ACB <= 1'b0; I916551CA30E7A94681BA2B3415BF85FA <= 1'b0; I4A3B5CD6A0CBD18332DCF8ECB309CC92
<= 1'b0; I2931854F66F4E6D5E96ED7D73266F38E <= 32'b0; IDA48F17DCE4BB1F6A04CBB23CCB4C3A5 <= {I15DA3B10E1E0658D2D01B744DF560903 {1'b0}};
IC93C4C87277AF77C73E35A77E14FC4B1 <= 1'b0; I54BE80AB8C90F3E5819921EF5354732A <= 1'b0; I7FA4C54BD6B551C794EE0EA588CBD4C7
<= 1'b0; I511F58CE0ACA83EE959D1BF6C4EAFA7F <= 1'b0; I623116EB4A13517E3733A1778B496560 <= 1'b0; I7E9516402D6933186513EB5B37336278
<= 8'b0; IA1EA4D4C05E159614ABC1E6D9CABE3BB <= 5'b0; I8916D921407646CE03BABA39B922EE09 <= 3'b0; I9C46AA186B65717669AB8B1F7ED02022
<= 1'b0; IE4E0DDAB16DD8E970672626428251866 <= 1'b0; IE12D7FB0707DA0B72DA8BD64B6FAEFEB <= 1'b0; I15C3BE43949B828A0A578329FE2EDE6B
<= 1'b0; IE655D625D2EB067AC17967E600BE5FBD <= 1'b0; IABBE7E409672B3D3CE209351AE63C530 <= 1'b0; I9962CDA8EE94C7BDFB23FE70815056E4
<= 1'b0; I7732946249B5963DFD9C95EC611A1D2C <= 1'b0; I54D7451A32675B2129629BC41778D6D6 <= 7'b0; I8AC99AB880823B01C00D137F89AABEF8
<= I3662C12143A4A1B904AC8798CEEF0125 ; I9B8138DCE156F7C31EB5914EF01F183C <= 1'b0; IB9A23596C80981B9B1CF7E12A76E71AC
<= 8'b0; I288715DFB3893A064D51571152559F12 <= 5'b0; I86B9557FA0123B8105E34300F4FCD447 <= 3'b0; I3EC90F87E70407C2A46DA25A8CA9065B
<= {IDE267FF256F75C9698907411CE334A5B {1'b0}}; I9E40C3A9F9E3CDFC05F95566701DFB02 <= 32'b0; ICFC6D424C8D5969FAC575FE0538F20F3
<= 1'b0; ICDFF33095CB0890DA2F167B63251EC67 <= 1'b0; IEDEC097EECBEE6B592219F6FEFFC7C2A <= 1'b0; I9E185DF5B08D79D1F56FD64627570AE0
<= 12'b0; I08AAFC572BC9A693B4E7C04DFD77FEAF <= 1'b0; I0C9005A5E5456704CE9C506A03373402 <= 8'b0; I5B0AA124C4ADA63A064AF2CAFA1098FD
<= {IDB9D60794264C5F8E5363941194A797B {1'b0}}; I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'b0; I83F18730E4735495B20E29C862E672F1
<= 64'b0; I18D210808E8E4FD4E19269D50B767EF6 <= 14'b0; I84B10D95B4B5E01F827E0D4D81BF476B <= 11'b0; I539C1D01FC349447001EB93E17D37611
<= 8'b0; I5B3BB6CF473F793585E2668A9A7136C8 <= 1'b0; I2C5E6805594DFF3B9EB915045ABF7575 <= 32'b0; I909A2BB1C99AC88EE130F2C2B36CD5AB
<= {I30AF2C9FF2EEDF02869CDAC1AAC433BC {1'b0}}; I893DF0D582AF0617B44879E65C202360 <= 1'b0; I2967174B668E2BB5A635A3F85DFF312B
<= 1'b0; I2212D954BC70C49C1F608E169DC873BC <= 1'b0; IC7779D4175ADF3F75C21392F9E824B6D <= {ID7C7F9F2E39BEBEE2ACFA8040034E48D {1'b0}};
IA6B00370F90E5BFE7B5D8852390CF107 <= 2'b0; I369C3845EEBC3367BADAF446789A185D <= 3'b0; I57E5F0C022683CA716D05ABE3408A469
<= 1'b0; IE7D8E2A0B7B7689804FFDF702BF724A6 <= 1'b0; I6F3C14B2AF4F4232F642DBEB36DCF09E <= 1'b0; I33F9C80AA280FFCBE2A2CB54C2056CC5
<= 1'b0; I5A4554E3FF0F3BAFC519CDF46237B987 <= {IDB9D60794264C5F8E5363941194A797B {1'b0}}; I074FD9C5AE408613B3750B75A6125486
<= 32'b0; IA934CBE3CC9AEBA0C32AA4C7EFA4954C <= 12'b0; I13C229A5BDE90D9F920D8F4D218106DE <= 4'b0; I037773E6A298229B4A19627ABA272E81
<= 1'b0; I0EBD58BCF1D55F648B20B722C25EA4A8 <= 1'b0; I30D7DB78C2B62A00872F044F1A2F39A2 <= {11{1'b0}}; I36FECBB048E15937DC767259CBABEDCB
<= 1'b0; end else begin I4A3B5CD6A0CBD18332DCF8ECB309CC92 <= IA886199C0F7609B072DAE171DFC98CD8 & I916551CA30E7A94681BA2B3415BF85FA ;
I2931854F66F4E6D5E96ED7D73266F38E <= I36824F33FF142FDE2AFE9BC4759DB690 ; I54BE80AB8C90F3E5819921EF5354732A <= I93AE636CE82DE94CB11ACCF59F8C2254 ;
I8AC99AB880823B01C00D137F89AABEF8 <= IF15E5692F18C2355720A228228564D0B ; I3EC90F87E70407C2A46DA25A8CA9065B <= I9F3623AEB414A15CECD2A8FD8791C79D ;
ICFC6D424C8D5969FAC575FE0538F20F3 <= IA886199C0F7609B072DAE171DFC98CD8 ; ICDFF33095CB0890DA2F167B63251EC67 <= (I3EC90F87E70407C2A46DA25A8CA9065B
>= I84B10D95B4B5E01F827E0D4D81BF476B ) ? ~I44B3CB0FFE4214C92C98CD6ECFC52D5A : 1'b0; I909A2BB1C99AC88EE130F2C2B36CD5AB
<= ICB518A59CAE27DDB6398AB22F5D74259 ; I893DF0D582AF0617B44879E65C202360 <= 1'b0; I2967174B668E2BB5A635A3F85DFF312B
<= (I909A2BB1C99AC88EE130F2C2B36CD5AB >= IA934CBE3CC9AEBA0C32AA4C7EFA4954C ) ? 1'b1 : 1'b0; I2212D954BC70C49C1F608E169DC873BC
<= 1'b0; I0EBD58BCF1D55F648B20B722C25EA4A8 <= 1'b0; if (IEDEC097EECBEE6B592219F6FEFFC7C2A == 1'b1) begin IEDEC097EECBEE6B592219F6FEFFC7C2A
<= (I9E185DF5B08D79D1F56FD64627570AE0 < 2) ? 1'b0 : IEDEC097EECBEE6B592219F6FEFFC7C2A ; I9E185DF5B08D79D1F56FD64627570AE0
<= (I9E185DF5B08D79D1F56FD64627570AE0 > 0) ? I9E185DF5B08D79D1F56FD64627570AE0 - 1 : {11{1'b0}}; I08AAFC572BC9A693B4E7C04DFD77FEAF
<= (I9E185DF5B08D79D1F56FD64627570AE0 < 2) ? 1'b1 : 1'b0; end if ((IEDEC097EECBEE6B592219F6FEFFC7C2A == 1'b1) &&
(IA886199C0F7609B072DAE171DFC98CD8 == 1'b0) && !((&I0C9005A5E5456704CE9C506A03373402 ) == 1'b1)) I0C9005A5E5456704CE9C506A03373402
<= I0C9005A5E5456704CE9C506A03373402 + 1; else if ((IEDEC097EECBEE6B592219F6FEFFC7C2A == 1'b0) && (IA886199C0F7609B072DAE171DFC98CD8
== 1'b1) && ((|I0C9005A5E5456704CE9C506A03373402 ) == 1'b1)) I0C9005A5E5456704CE9C506A03373402 <= I0C9005A5E5456704CE9C506A03373402
- 1; if (IA886199C0F7609B072DAE171DFC98CD8 == 1'b1) I9E40C3A9F9E3CDFC05F95566701DFB02 <= I36824F33FF142FDE2AFE9BC4759DB690 ;
case (I8AC99AB880823B01C00D137F89AABEF8 ) I3662C12143A4A1B904AC8798CEEF0125 : begin I916551CA30E7A94681BA2B3415BF85FA
<= 1'b0; if (I9F3623AEB414A15CECD2A8FD8791C79D > 2) begin I08AAFC572BC9A693B4E7C04DFD77FEAF <= 1'b0; I9E185DF5B08D79D1F56FD64627570AE0
<= 11'h003; IEDEC097EECBEE6B592219F6FEFFC7C2A <= 1'b1; end end I257DF24B77C5CA85F676E7FFA065CE94 : begin IDA48F17DCE4BB1F6A04CBB23CCB4C3A5
<= I15DA3B10E1E0658D2D01B744DF560903 - 1; I83F18730E4735495B20E29C862E672F1 <= {64{1'b0}}; I893DF0D582AF0617B44879E65C202360
<= 1'b0; end I54DD54FD7FB944705CE08C2B291B87A7 : begin I7FA4C54BD6B551C794EE0EA588CBD4C7 <= 1'b0; I511F58CE0ACA83EE959D1BF6C4EAFA7F
<= I9E40C3A9F9E3CDFC05F95566701DFB02 [30]; I623116EB4A13517E3733A1778B496560 <= ~I9E40C3A9F9E3CDFC05F95566701DFB02 [29];
IEDEC097EECBEE6B592219F6FEFFC7C2A <= I9E40C3A9F9E3CDFC05F95566701DFB02 [29]; I18D210808E8E4FD4E19269D50B767EF6 <=
I9E40C3A9F9E3CDFC05F95566701DFB02 [23:10]; I84B10D95B4B5E01F827E0D4D81BF476B <= {1'b0, I9E40C3A9F9E3CDFC05F95566701DFB02 [10:0]};
I9C46AA186B65717669AB8B1F7ED02022 <= ((I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I81D26620360085DCC2783D5734873451 )
|| (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == IA3187A41E33086C9DA805D8C67004992 )) ? 1'b1 : 1'b0; IE4E0DDAB16DD8E970672626428251866
<= ((I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I2C8281C2456BAC869C04372CE6A7C50E ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24]
== I8CD6057CFBD7215340EF60C41A0C63EC )) ? 1'b1 : 1'b0; IE12D7FB0707DA0B72DA8BD64B6FAEFEB <= ((I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24]
== I6A62FD6104E281B8714322DB8CCB5FE3 ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I85B0192F2AC4464C88E2C93352FE6696 )
|| (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I78DDE5821936F928E302A8BA3C3138EE ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24]
== I41F249A62806D544C38454CA2D10750D )) ? 1'b1 : 1'b0; I15C3BE43949B828A0A578329FE2EDE6B <= ((I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24]
== I34EF8B0D0058C1876C19361DBBAC62DC ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == IB83A8F7EA6693A633C486F9CA18003BB ))
? 1'b1 : 1'b0; IE655D625D2EB067AC17967E600BE5FBD <= ((I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I8F0EB88EC813DC0B3105F31BABD34B79 )
|| (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I877B2A234FC10EC8A4A2F0A90F6EAE6C ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24]
== IEC10F95DD42CAF869EFB03BDF59BE8EB ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I2E664E814B6AA2CBCE57FBCE2A354435 ))
? 1'b1 : 1'b0; IABBE7E409672B3D3CE209351AE63C530 <= (((I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] & 8'hf0) == IBC983AF54FD90EA2AA9E3DD139A3B818 )
|| ((I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] & 8'hf0) == I361F321AEF89DD0EF2CEAC65B8B042D8 )) ? 1'b1 : 1'b0; I9962CDA8EE94C7BDFB23FE70815056E4
<= ((I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I8F0EB88EC813DC0B3105F31BABD34B79 ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24]
== I877B2A234FC10EC8A4A2F0A90F6EAE6C ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I81D26620360085DCC2783D5734873451 )
|| (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == IA3187A41E33086C9DA805D8C67004992 ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24]
== I2C8281C2456BAC869C04372CE6A7C50E ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I8CD6057CFBD7215340EF60C41A0C63EC )
|| (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I34EF8B0D0058C1876C19361DBBAC62DC ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24]
== IB83A8F7EA6693A633C486F9CA18003BB )) ? 1'b1 : 1'b0; if (I9E40C3A9F9E3CDFC05F95566701DFB02 [29]) begin I08AAFC572BC9A693B4E7C04DFD77FEAF
<= 1'b0; I9E185DF5B08D79D1F56FD64627570AE0 <= 11'h001; IEDEC097EECBEE6B592219F6FEFFC7C2A <= 1'b1; end end I962A83F6AB78F0114DD9D85409B29E8F
: begin I11FD35FED78BCB8861FACB9A1E3A4C35 <= I9E40C3A9F9E3CDFC05F95566701DFB02 [3:0]; IC52F3B77F7E45A74323561D6A6F6028A
<= I9E40C3A9F9E3CDFC05F95566701DFB02 [7:4]; I539C1D01FC349447001EB93E17D37611 <= I9E40C3A9F9E3CDFC05F95566701DFB02 [15:8];
IB9A23596C80981B9B1CF7E12A76E71AC <= I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24]; I288715DFB3893A064D51571152559F12
<= I9E40C3A9F9E3CDFC05F95566701DFB02 [23:19]; I86B9557FA0123B8105E34300F4FCD447 <= I9E40C3A9F9E3CDFC05F95566701DFB02 [18:16];
I30D7DB78C2B62A00872F044F1A2F39A2 <= {((I84B10D95B4B5E01F827E0D4D81BF476B [9:0] == 0) ? 1'b1 : 1'b0), I84B10D95B4B5E01F827E0D4D81BF476B [9:0]};
I84B10D95B4B5E01F827E0D4D81BF476B [10] <= (I84B10D95B4B5E01F827E0D4D81BF476B [9:0] == 0) ? 1'b1 : 1'b0; end IA4997CC969740D4CF1FC8E4E9C2B5DA7
: begin I71DBDE411F9CED520FD43A4EF5CBD656 <= (I84B10D95B4B5E01F827E0D4D81BF476B [1:0] == 2'b00) ? I84B10D95B4B5E01F827E0D4D81BF476B [10:2]
: I84B10D95B4B5E01F827E0D4D81BF476B [10:2] + 1; I7E9516402D6933186513EB5B37336278 <= I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24];
IA1EA4D4C05E159614ABC1E6D9CABE3BB <= I9E40C3A9F9E3CDFC05F95566701DFB02 [23:19]; I8916D921407646CE03BABA39B922EE09
<= I9E40C3A9F9E3CDFC05F95566701DFB02 [18:16]; IC7779D4175ADF3F75C21392F9E824B6D <= {ID7C7F9F2E39BEBEE2ACFA8040034E48D {1'b0}};
IA934CBE3CC9AEBA0C32AA4C7EFA4954C <= I30D7DB78C2B62A00872F044F1A2F39A2 ; if (I9C46AA186B65717669AB8B1F7ED02022 |
IE4E0DDAB16DD8E970672626428251866 ) begin I83F18730E4735495B20E29C862E672F1 [31:0] <= {17'b0, I9E40C3A9F9E3CDFC05F95566701DFB02 [18:16],
I9E40C3A9F9E3CDFC05F95566701DFB02 [11:0]}; I83F18730E4735495B20E29C862E672F1 [63:32] <= {32{1'b0}}; end else begin
I83F18730E4735495B20E29C862E672F1 [31:0] <= I9E40C3A9F9E3CDFC05F95566701DFB02 ; I83F18730E4735495B20E29C862E672F1 [63:32]
<= {32{1'b0}}; end case (IC52F3B77F7E45A74323561D6A6F6028A ) 4'b0100, 4'b0101, 4'b0110, 4'b0111 : case (I11FD35FED78BCB8861FACB9A1E3A4C35 )
4'b0010, 4'b0110, 4'b1010, 4'b1110 : I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd2; 4'b0100, 4'b1100 : I93F6D99D18FD6FF40EF5AD5288D5C88E
<= 4'd3; 4'b1000 : I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd4; default I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd1;
endcase 4'b0010, 4'b0011 : case (I11FD35FED78BCB8861FACB9A1E3A4C35 ) 4'b0010, 4'b0110, 4'b1010, 4'b1110 : I93F6D99D18FD6FF40EF5AD5288D5C88E
<= 4'd3; 4'b0100, 4'b1100 : I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd4; 4'b1000 : I93F6D99D18FD6FF40EF5AD5288D5C88E
<= 4'd5; default I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd2; endcase 4'b0001 : case (I11FD35FED78BCB8861FACB9A1E3A4C35 )
4'b0010, 4'b0110, 4'b1010, 4'b1110 : I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd4; 4'b0100, 4'b1100 : I93F6D99D18FD6FF40EF5AD5288D5C88E
<= 4'd5; 4'b1000 : I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd6; default I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd3;
endcase 4'b0000 : case (I11FD35FED78BCB8861FACB9A1E3A4C35 ) 4'b0000, 4'b0001, 4'b0010, 4'b0100, 4'b1000 : I93F6D99D18FD6FF40EF5AD5288D5C88E
<= 4'd3; 4'b0011, 4'b0110, 4'b1100 : I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd2; 4'b0101, 4'b0111, 4'b1010, 4'b1110
: I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd1; default I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd0; endcase default
case (I11FD35FED78BCB8861FACB9A1E3A4C35 ) 4'b0010, 4'b0110, 4'b1010, 4'b1110 : I93F6D99D18FD6FF40EF5AD5288D5C88E
<= 4'd1; 4'b0100, 4'b1100 : I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd2; 4'b1000 : I93F6D99D18FD6FF40EF5AD5288D5C88E
<= 4'd3; default I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd0; endcase endcase end I8EBFD17705709FF6F2CAA85EA87D66D4
: begin if (ICFC6D424C8D5969FAC575FE0538F20F3 ) I83F18730E4735495B20E29C862E672F1 <= {I83F18730E4735495B20E29C862E672F1 [31:0],
I9E40C3A9F9E3CDFC05F95566701DFB02 }; end I56AC73D28E70D2F78200164359CC0E9A : begin I0FF03F7D70F3047C91A55F9744DDD7AE
<= (IB9A23596C80981B9B1CF7E12A76E71AC == IFF5E23C5A17BB678C108274E28C56424 ) ? 1'b1 : 1'b0; IC93C4C87277AF77C73E35A77E14FC4B1
<= (I288715DFB3893A064D51571152559F12 == IDE425A12275C43D9056DCF647A2D8258 ) ? 1'b1 : 1'b0; if (IDA48F17DCE4BB1F6A04CBB23CCB4C3A5 )
IDA48F17DCE4BB1F6A04CBB23CCB4C3A5 <= IDA48F17DCE4BB1F6A04CBB23CCB4C3A5 - 1; end I499DB4E92AEE1C97FE024F6FD8CDEB8A
: begin IAC85A6B0EE1F3079B60C115CB476DF06 <= {I30D7DB78C2B62A00872F044F1A2F39A2 [9:0], 2'b00} - I93F6D99D18FD6FF40EF5AD5288D5C88E ;
I916551CA30E7A94681BA2B3415BF85FA <= IE12D7FB0707DA0B72DA8BD64B6FAEFEB & ((I7E9516402D6933186513EB5B37336278 ==
IFF5E23C5A17BB678C108274E28C56424 ) ? 1'b1 : 1'b0) & ((IA1EA4D4C05E159614ABC1E6D9CABE3BB == IDE425A12275C43D9056DCF647A2D8258 )
? 1'b1 : 1'b0); I7732946249B5963DFD9C95EC611A1D2C <= ~I93FEA934E2F91A4D5E773376B9B26FED ; I5B0AA124C4ADA63A064AF2CAFA1098FD
<= (IE655D625D2EB067AC17967E600BE5FBD | I15C3BE43949B828A0A578329FE2EDE6B ) ? I7E600D684E83043922C1FE27CC6213E4
: {IDB9D60794264C5F8E5363941194A797B {1'b0}}; end IABEE3580E02F366EC5560A9CFC5CC953 : begin if (ICDFF33095CB0890DA2F167B63251EC67
== 1'b1) begin I08AAFC572BC9A693B4E7C04DFD77FEAF <= 1'b0; I9E185DF5B08D79D1F56FD64627570AE0 <= I84B10D95B4B5E01F827E0D4D81BF476B ;
IEDEC097EECBEE6B592219F6FEFFC7C2A <= 1'b1; end end I174E152AA0198C30C57B401C947D37C1 : begin IA6B00370F90E5BFE7B5D8852390CF107
<= I6768A159F7F57847F9535CB8B8B382D8 ; I57E5F0C022683CA716D05ABE3408A469 <= I9C46AA186B65717669AB8B1F7ED02022 ;
IE7D8E2A0B7B7689804FFDF702BF724A6 <= IE4E0DDAB16DD8E970672626428251866 ; I6F3C14B2AF4F4232F642DBEB36DCF09E <= IE12D7FB0707DA0B72DA8BD64B6FAEFEB ;
I369C3845EEBC3367BADAF446789A185D <= (I84B10D95B4B5E01F827E0D4D81BF476B == 1) ? IEE94C2462F89091D3C62992327532D1E
: I88A97019335E3F57955B11E67DFFCD65 ; I33F9C80AA280FFCBE2A2CB54C2056CC5 <= IABBE7E409672B3D3CE209351AE63C530 ; I5A4554E3FF0F3BAFC519CDF46237B987
<= I5B0AA124C4ADA63A064AF2CAFA1098FD ; I074FD9C5AE408613B3750B75A6125486 <= (I511F58CE0ACA83EE959D1BF6C4EAFA7F ==
1'b1) ? I36824F33FF142FDE2AFE9BC4759DB690 : 32'b0; I13C229A5BDE90D9F920D8F4D218106DE <= I11FD35FED78BCB8861FACB9A1E3A4C35 ;
I037773E6A298229B4A19627ABA272E81 <= ((IA886199C0F7609B072DAE171DFC98CD8 == 1'b1) || (I511F58CE0ACA83EE959D1BF6C4EAFA7F
== 1'b0)) ? 1'b1 : 1'b0; I0EBD58BCF1D55F648B20B722C25EA4A8 <= 1'b1; I36FECBB048E15937DC767259CBABEDCB <= I511F58CE0ACA83EE959D1BF6C4EAFA7F ;
if (IE12D7FB0707DA0B72DA8BD64B6FAEFEB ) IC7779D4175ADF3F75C21392F9E824B6D [14:0] <= {I86B9557FA0123B8105E34300F4FCD447 ,
I83F18730E4735495B20E29C862E672F1 [11:2], 2'b00}; else IC7779D4175ADF3F75C21392F9E824B6D <= {I83F18730E4735495B20E29C862E672F1 [ID7C7F9F2E39BEBEE2ACFA8040034E48D
- 1:2], 2'b00}; end I3C15F904BACDB851EFC4C548820E98B8 : begin I2212D954BC70C49C1F608E169DC873BC <= I07B0EBE8FBC21BDBE894D73C90EDC5AB ;
if (I07B0EBE8FBC21BDBE894D73C90EDC5AB ) begin I893DF0D582AF0617B44879E65C202360 <= (I369C3845EEBC3367BADAF446789A185D
== IEE94C2462F89091D3C62992327532D1E ) ? 1'b1 : 1'b0; I369C3845EEBC3367BADAF446789A185D <= (IA934CBE3CC9AEBA0C32AA4C7EFA4954C
== 2) ? IEE94C2462F89091D3C62992327532D1E : I88A97019335E3F57955B11E67DFFCD65 ; I13C229A5BDE90D9F920D8F4D218106DE
<= 4'b1111; IA934CBE3CC9AEBA0C32AA4C7EFA4954C <= IA934CBE3CC9AEBA0C32AA4C7EFA4954C - 1; if (I9B8138DCE156F7C31EB5914EF01F183C )
I2C5E6805594DFF3B9EB915045ABF7575 <= I44109A75F9883AA09218902DA5B2CBB3 ; else I2C5E6805594DFF3B9EB915045ABF7575
<= {32{1'b1}}; if (I369C3845EEBC3367BADAF446789A185D == IEE94C2462F89091D3C62992327532D1E ) begin IC7779D4175ADF3F75C21392F9E824B6D
<= {ID7C7F9F2E39BEBEE2ACFA8040034E48D {1'b0}}; I074FD9C5AE408613B3750B75A6125486 <= 32'b0; IA6B00370F90E5BFE7B5D8852390CF107
<= 2'b0; I369C3845EEBC3367BADAF446789A185D <= 3'b0; I57E5F0C022683CA716D05ABE3408A469 <= 1'b0; IE7D8E2A0B7B7689804FFDF702BF724A6
<= 1'b0; I6F3C14B2AF4F4232F642DBEB36DCF09E <= 1'b0; I33F9C80AA280FFCBE2A2CB54C2056CC5 <= 1'b0; I5A4554E3FF0F3BAFC519CDF46237B987
<= {IDB9D60794264C5F8E5363941194A797B {1'b0}}; I13C229A5BDE90D9F920D8F4D218106DE <= 4'b0; I037773E6A298229B4A19627ABA272E81
<= 1'b0; I36FECBB048E15937DC767259CBABEDCB <= 1'b0; end end end I29C10DD8DAC8AB31273614BA27A5E29C : begin if (I07B0EBE8FBC21BDBE894D73C90EDC5AB )
begin I369C3845EEBC3367BADAF446789A185D <= (IA934CBE3CC9AEBA0C32AA4C7EFA4954C == 2) ? IEE94C2462F89091D3C62992327532D1E
: I88A97019335E3F57955B11E67DFFCD65 ; I13C229A5BDE90D9F920D8F4D218106DE <= (IA934CBE3CC9AEBA0C32AA4C7EFA4954C ==
2) ? IC52F3B77F7E45A74323561D6A6F6028A : 4'b1111; IA934CBE3CC9AEBA0C32AA4C7EFA4954C <= IA934CBE3CC9AEBA0C32AA4C7EFA4954C
- 1; if (I369C3845EEBC3367BADAF446789A185D == IEE94C2462F89091D3C62992327532D1E ) begin IC7779D4175ADF3F75C21392F9E824B6D
<= {ID7C7F9F2E39BEBEE2ACFA8040034E48D {1'b0}}; I074FD9C5AE408613B3750B75A6125486 <= 32'b0; IA6B00370F90E5BFE7B5D8852390CF107
<= 2'b0; I369C3845EEBC3367BADAF446789A185D <= 3'b0; I57E5F0C022683CA716D05ABE3408A469 <= 1'b0; IE7D8E2A0B7B7689804FFDF702BF724A6
<= 1'b0; I6F3C14B2AF4F4232F642DBEB36DCF09E <= 1'b0; I33F9C80AA280FFCBE2A2CB54C2056CC5 <= 1'b0; I5A4554E3FF0F3BAFC519CDF46237B987
<= {IDB9D60794264C5F8E5363941194A797B {1'b0}}; I074FD9C5AE408613B3750B75A6125486 <= 32'b0; I13C229A5BDE90D9F920D8F4D218106DE
<= 4'b0; I037773E6A298229B4A19627ABA272E81 <= 1'b0; I36FECBB048E15937DC767259CBABEDCB <= 1'b0; end else begin I074FD9C5AE408613B3750B75A6125486
<= I36824F33FF142FDE2AFE9BC4759DB690 ; end end end IF5A7A7CE92502E2DF9F0601605A38637 : begin if (I9962CDA8EE94C7BDFB23FE70815056E4 )
begin if (~IA85D446CD214F6B3CE6418205432D870 ) I26F46DF735C89C3DA76F7F404A5F650F <= 1'b1; if (I511F58CE0ACA83EE959D1BF6C4EAFA7F
& ~I69B8FD7561F9CA8AAF4E50C5B2DCF850 ) begin IBFF7FD594C616C9EBAD12448149DA576 <= I71DBDE411F9CED520FD43A4EF5CBD656 ;
I0C9CC98CD774EDC9DF9AB513E5A8FB57 <= 1'b1; end end else if (~IE12D7FB0707DA0B72DA8BD64B6FAEFEB ) begin if (~I45A8F29589769D54C9D702481065CB45 )
IF9A51F60DF053D68A5D57FECB5AB7ACB <= 1'b1; if (I511F58CE0ACA83EE959D1BF6C4EAFA7F & ~IBB8FE5B389C0BD7BA64F2E05FCDC4485 )begin
I5AF6C20F3950D58007B9C0BEA7C87198 <= I71DBDE411F9CED520FD43A4EF5CBD656 ; I533559C7D3A6FC7D4A2E49A02AFC9137 <= 1'b1;
end end if (I50AC25E9687F891BB7188EED025C1323 ) if ((I623116EB4A13517E3733A1778B496560 && (!I511F58CE0ACA83EE959D1BF6C4EAFA7F
|| (I511F58CE0ACA83EE959D1BF6C4EAFA7F && ~I84B10D95B4B5E01F827E0D4D81BF476B [0]))) || (!I623116EB4A13517E3733A1778B496560
&& I511F58CE0ACA83EE959D1BF6C4EAFA7F && I84B10D95B4B5E01F827E0D4D81BF476B [0])) begin I08AAFC572BC9A693B4E7C04DFD77FEAF
<= 1'b0; I9E185DF5B08D79D1F56FD64627570AE0 <= 11'h001; IEDEC097EECBEE6B592219F6FEFFC7C2A <= 1'b1; end end I5021A214EB457E909E76C621F6DD12B1
: begin IBFF7FD594C616C9EBAD12448149DA576 <= 8'b0; I0C9CC98CD774EDC9DF9AB513E5A8FB57 <= 1'b0; I26F46DF735C89C3DA76F7F404A5F650F
<= 1'b0; I5AF6C20F3950D58007B9C0BEA7C87198 <= 8'b0; I533559C7D3A6FC7D4A2E49A02AFC9137 <= 1'b0; IF9A51F60DF053D68A5D57FECB5AB7ACB
<= 1'b0; end I05E305FFF5B6CDE122F8935EE521D523 : begin I5B3BB6CF473F793585E2668A9A7136C8 <= ~I5B3BB6CF473F793585E2668A9A7136C8
| (I5B3BB6CF473F793585E2668A9A7136C8 & ~I9F4F7E2C4A4A8FB2780021EDF6E4ADEF ); end IFAC7B411ECB5421590DDAA0B7B34F238
: begin if (I511F58CE0ACA83EE959D1BF6C4EAFA7F ) if (ICDFF33095CB0890DA2F167B63251EC67 ) begin I08AAFC572BC9A693B4E7C04DFD77FEAF
<= 1'b0; I9E185DF5B08D79D1F56FD64627570AE0 <= I84B10D95B4B5E01F827E0D4D81BF476B ; IEDEC097EECBEE6B592219F6FEFFC7C2A
<= 1'b1; end end I6EA1237B063AFA6C82E354D0001BEF41 : begin I7FA4C54BD6B551C794EE0EA588CBD4C7 <= 1'b1; I9B8138DCE156F7C31EB5914EF01F183C
<= I9119CE851F731CBC5834D0370CCA6908 [I6345C4C803C15670FB2665AEA7AA4E33 ] | I9C46AA186B65717669AB8B1F7ED02022 ;
if (I511F58CE0ACA83EE959D1BF6C4EAFA7F | I7732946249B5963DFD9C95EC611A1D2C ) I2C5E6805594DFF3B9EB915045ABF7575 <=
{I6A62FD6104E281B8714322DB8CCB5FE3 , I18D210808E8E4FD4E19269D50B767EF6 , 10'b0}; else if (IE655D625D2EB067AC17967E600BE5FBD )
I2C5E6805594DFF3B9EB915045ABF7575 <= {I85B0192F2AC4464C88E2C93352FE6696 , I18D210808E8E4FD4E19269D50B767EF6 , I30D7DB78C2B62A00872F044F1A2F39A2 [9:0]};
else I2C5E6805594DFF3B9EB915045ABF7575 <= {I85B0192F2AC4464C88E2C93352FE6696 , I18D210808E8E4FD4E19269D50B767EF6 ,
10'b01}; I2212D954BC70C49C1F608E169DC873BC <= 1'b1; case (I11FD35FED78BCB8861FACB9A1E3A4C35 ) 4'b0010, 4'b0110,
4'b1010, 4'b1110 : I54D7451A32675B2129629BC41778D6D6 <= {I83F18730E4735495B20E29C862E672F1 [6:2], 2'b01}; 4'b0100,
4'b1100 : I54D7451A32675B2129629BC41778D6D6 <= {I83F18730E4735495B20E29C862E672F1 [6:2], 2'b10}; 4'b1000 : I54D7451A32675B2129629BC41778D6D6
<= {I83F18730E4735495B20E29C862E672F1 [6:2], 2'b11}; default I54D7451A32675B2129629BC41778D6D6 <= I83F18730E4735495B20E29C862E672F1 [6:0];
endcase end ID1D4A1F29119D84947D94DCCD5BDF6A9 : begin if (I7732946249B5963DFD9C95EC611A1D2C ) if (IE655D625D2EB067AC17967E600BE5FBD )
I2C5E6805594DFF3B9EB915045ABF7575 <= {IC4C940842A3072C3A9C40616C6A213F2 , IE8010EDEC4159FBD688A550900D0006D , I6345C4C803C15670FB2665AEA7AA4E33 ,
ID2A58EC9E1C805C9EA9CF0D05ACFD523 , 1'b0, IAC85A6B0EE1F3079B60C115CB476DF06 }; else I2C5E6805594DFF3B9EB915045ABF7575
<= {IC4C940842A3072C3A9C40616C6A213F2 , IE8010EDEC4159FBD688A550900D0006D , I6345C4C803C15670FB2665AEA7AA4E33 ,
ID2A58EC9E1C805C9EA9CF0D05ACFD523 , 1'b0, 12'h004}; else if (IE655D625D2EB067AC17967E600BE5FBD ) I2C5E6805594DFF3B9EB915045ABF7575
<= {IC4C940842A3072C3A9C40616C6A213F2 , IE8010EDEC4159FBD688A550900D0006D , I6345C4C803C15670FB2665AEA7AA4E33 ,
IF79BEED009A88E1D471FE1CEC77A7604 , 1'b0, IAC85A6B0EE1F3079B60C115CB476DF06 }; else I2C5E6805594DFF3B9EB915045ABF7575
<= {IC4C940842A3072C3A9C40616C6A213F2 , IE8010EDEC4159FBD688A550900D0006D , I6345C4C803C15670FB2665AEA7AA4E33 ,
IF79BEED009A88E1D471FE1CEC77A7604 , 1'b0, 12'h004}; I2212D954BC70C49C1F608E169DC873BC <= 1'b1; end IF86E23BE5E6D56399363666A2BDC7A6A
: begin if (IE655D625D2EB067AC17967E600BE5FBD ) I2C5E6805594DFF3B9EB915045ABF7575 <= {IB9A23596C80981B9B1CF7E12A76E71AC ,
I288715DFB3893A064D51571152559F12 , I86B9557FA0123B8105E34300F4FCD447 , I539C1D01FC349447001EB93E17D37611 , 1'b0,
I54D7451A32675B2129629BC41778D6D6 }; else I2C5E6805594DFF3B9EB915045ABF7575 <= {IB9A23596C80981B9B1CF7E12A76E71AC ,
I288715DFB3893A064D51571152559F12 , I86B9557FA0123B8105E34300F4FCD447 , I539C1D01FC349447001EB93E17D37611 , 1'b0,
7'b0}; I893DF0D582AF0617B44879E65C202360 <= I7732946249B5963DFD9C95EC611A1D2C | I511F58CE0ACA83EE959D1BF6C4EAFA7F ;
I2212D954BC70C49C1F608E169DC873BC <= 1'b1; end I264B836E51E7F23F603A59DFDC8D2C8A : begin I2C5E6805594DFF3B9EB915045ABF7575
<= 32'b0; I893DF0D582AF0617B44879E65C202360 <= 1'b0; I2212D954BC70C49C1F608E169DC873BC <= 1'b0; end endcase end
end endmodule 
  module I1F8444FEC9FE4C651C698EE6099B529D #( parameter IB71844FFA3AB85FEF45EAB4D35395752 = 256, parameter IDB9D60794264C5F8E5363941194A797B
= 3, parameter ID7C7F9F2E39BEBEE2ACFA8040034E48D = 16 ) ( input wire ICCFB0F435B37370076102F325BC08D20 , input wire
I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire I69B8FD7561F9CA8AAF4E50C5B2DCF850 , input wire IA85D446CD214F6B3CE6418205432D870 ,
input wire IBB8FE5B389C0BD7BA64F2E05FCDC4485 , input wire I45A8F29589769D54C9D702481065CB45 , input wire [7:0] IFF5E23C5A17BB678C108274E28C56424 ,
input wire [4:0] IDE425A12275C43D9056DCF647A2D8258 , input wire [2:0] I65B14714ECFCC218D3A788DF7696216B , input
wire [2:0] IA1F0CBEC8E9EAD83D0098DD96A1EFC32 , input wire IFC18758E8987A9913FD94A5DFEE774E2 , input wire IF5E7E4E58741BF3FE58442AB377ED57F ,
input wire IF5B4924BEAEA6935367AC2739021882F , input wire I7985A5A43CBBBC8E0D3FCFEE38DDF221 , input wire [IDB9D60794264C5F8E5363941194A797B
- 1:0] I7E600D684E83043922C1FE27CC6213E4 , input wire I93AE636CE82DE94CB11ACCF59F8C2254 , input wire [7:0] I9119CE851F731CBC5834D0370CCA6908 ,
input wire [$clog2(IB71844FFA3AB85FEF45EAB4D35395752 + 1) - 1:0] I9F3623AEB414A15CECD2A8FD8791C79D , input wire
[63:0] I36824F33FF142FDE2AFE9BC4759DB690 , input wire I5E84ED10AD623502BC750C5E797D1428 , input wire IA886199C0F7609B072DAE171DFC98CD8 ,
input wire IA067043029572C8598E352E0A66EA337 , input wire [$clog2(IB71844FFA3AB85FEF45EAB4D35395752 + 1) - 1:0]
ICB518A59CAE27DDB6398AB22F5D74259 , input wire I9F4F7E2C4A4A8FB2780021EDF6E4ADEF , input wire I07B0EBE8FBC21BDBE894D73C90EDC5AB ,
input wire I44B3CB0FFE4214C92C98CD6ECFC52D5A , input wire [63:0] I3D6C771D05CA1A769E61302C086494B8 , output wire
[7:0] IC2E260CA356C994048CCB108C7E359D1 , output wire [7:0] IE707B5D4A74BA1BD745B52E0C07932C0 , output wire I6E70C748D9C56227AB1182F36658AE5C ,
output wire I59B23598E8ADE1982F184EF67BEB0979 , output wire I33E409903692F5ECA2EC3553F9D1659E , output wire I437E57D42FB91B674CCBCC915BF9D653 ,
output wire I55AFDDE17B53D7F65849D39B02B07417 , output wire [63:0] I65FE2DB4E1CB5A488A45D60041AB5F64 , output wire
[63:0] I0C796C206FE7060B578156D0110461EB , output wire IFC86A6522A8CA080A0DB7F384D9CE6FA , output wire I484F77D7967D25736EB27A0ED76CCB5F ,
output wire I7E0431D7F1A92C0ED1F030F36BF809B7 , output wire I3E6965EC606FD6C2871F2C0993204C57 , output wire IFF25B820DFD457D71B32B130ABE5DA3F ,
output wire I20FA57C9A87CB2AA26088D9FA1743F70 , output wire I51C881E8B9B36D7A724BC7B8EC533957 , output wire [7:0]
ID3E7F4B58943229FEE6313A36B3F8693 , output wire [4:0] I1FDEC1735547330C00A0B8DFE1FB10C3 , output wire [2:0] IBD6A65D48B4A68CA0D2A82F79053757B ,
output wire I15EC78E3DE1101BFF2B227962683E113 , output wire [63:0] I7C4DADE2C05F6DCECCAF7AD6F7BF2FF8 , output wire
IEEFA85D6664F09687B5CA591C701DC34 , output wire ID4A284C76C6EABEEBA8E0AE18003FBAC , output wire I6010C20131B976554A498745FEEEB580 ,
output wire [ID7C7F9F2E39BEBEE2ACFA8040034E48D - 1:0] I46E8CA15DC1E8B3B2200999A53029704 , output wire [1:0] IEC45B60C7D1A49FFA84D3F5D121A2579 ,
output wire [2:0] I9AF46E2AA924FA7E0F5D7290324BABF9 , output wire I59D9A9A677978229C1F87AA1A3A0C304 , output wire
I9301CE4E9B877D08EDBD1584D6BE017A , output wire I51698892CBD372EE66AF3EA4D0ECE23F , output wire I1347408C9E757F34EA4D78F53447BD9B ,
output wire [IDB9D60794264C5F8E5363941194A797B - 1:0] I2BE88607F3C31B47400F3A35E08B7EAD , output wire [63:0] I7D901091F9E0741061C75B54467D48A0 ,
output wire I7AEBDB3D2CD4891A528BA81F5F54B20D , output wire [10:0] ID16819FEAA95700005E383E7DA0C8E13 , output wire
[3:0] IE0337CA803FBA20F38A0CD2A900C6534 , output wire [3:0] I592A6A3BA99B09C24695C7A609F9053F , output wire [3:0]
I40EF39BB4F4F4A031C8FD1026EF53063 , output wire I42427E866FF31BC28E35C71EC172E26B , output wire I368749E68EAF9F462385FAD36180A9FE
); `include "pcisig_constants.v"
`include "wishbone_utils.v"
 localparam I15DA3B10E1E0658D2D01B744DF560903 = 3; localparam I1797388B2E6E3CB5EE600DD85605F982 = $clog2(I15DA3B10E1E0658D2D01B744DF560903 );
localparam I63F1EFA9086319A16127622F3CE8B7D0 = $clog2(IB71844FFA3AB85FEF45EAB4D35395752 + 1); localparam I3662C12143A4A1B904AC8798CEEF0125
= 5'b00000, I257DF24B77C5CA85F676E7FFA065CE94 = 5'b00001, I67E645B7D6135C108074CF368E9BB834 = 5'b00010, IFE893DBF9067A0DA39E179005AD783C4
= 5'b00011, I56AC73D28E70D2F78200164359CC0E9A = 5'b00100, I499DB4E92AEE1C97FE024F6FD8CDEB8A = 5'b00101, IABEE3580E02F366EC5560A9CFC5CC953
= 5'b00110, I2D358EAE916810B434B6C76F7C7C5673 = 5'b00111, I174E152AA0198C30C57B401C947D37C1 = 5'b01000, I3C15F904BACDB851EFC4C548820E98B8
= 5'b01001, I61A7D75570E89738696B9598A883C1CD = 5'b01010, I29C10DD8DAC8AB31273614BA27A5E29C = 5'b01011, IF5A7A7CE92502E2DF9F0601605A38637
= 5'b01100, I5021A214EB457E909E76C621F6DD12B1 = 5'b01101, IFAC7B411ECB5421590DDAA0B7B34F238 = 5'b01110, I248DCDE6260EE21AB43E9E1EF6D603EF
= 5'b01111, IC495D10CCC7452A18D769BDD99794652 = 5'b10000, IEAE55E29AC7D8EC5093BF4C91D5CFFCE = 5'b10001, I6EA1237B063AFA6C82E354D0001BEF41
= 5'b10010, I070181DB2ED3EDD3633DB4E93B8E42A5 = 5'b10011, I2263EE3B1CDD9957F685B729A9639643 = 5'b10100, I05E305FFF5B6CDE122F8935EE521D523
= 5'b10101;  reg [3:0] I11FD35FED78BCB8861FACB9A1E3A4C35 ; reg [3:0] IC52F3B77F7E45A74323561D6A6F6028A ; reg I0FF03F7D70F3047C91A55F9744DDD7AE ;
reg [11:0] IAC85A6B0EE1F3079B60C115CB476DF06 ; reg [8:0] I71DBDE411F9CED520FD43A4EF5CBD656 ; reg [7:0] IBFF7FD594C616C9EBAD12448149DA576 ;
reg I0C9CC98CD774EDC9DF9AB513E5A8FB57 ; reg I26F46DF735C89C3DA76F7F404A5F650F ; reg [7:0] I5AF6C20F3950D58007B9C0BEA7C87198 ;
reg I533559C7D3A6FC7D4A2E49A02AFC9137 ; reg IF9A51F60DF053D68A5D57FECB5AB7ACB ; reg I916551CA30E7A94681BA2B3415BF85FA ;
reg I4A3B5CD6A0CBD18332DCF8ECB309CC92 ; reg [63:0] I2931854F66F4E6D5E96ED7D73266F38E ; reg [I1797388B2E6E3CB5EE600DD85605F982
- 1:0] IDA48F17DCE4BB1F6A04CBB23CCB4C3A5 ; reg IC93C4C87277AF77C73E35A77E14FC4B1 ; reg I54BE80AB8C90F3E5819921EF5354732A ;
reg IF4B2F356412545C21578876129150C2F ; reg I511F58CE0ACA83EE959D1BF6C4EAFA7F ; reg [7:0] I7E9516402D6933186513EB5B37336278 ;
reg [4:0] IA1EA4D4C05E159614ABC1E6D9CABE3BB ; reg [2:0] I8916D921407646CE03BABA39B922EE09 ; reg I7FA4C54BD6B551C794EE0EA588CBD4C7 ;
reg I9C46AA186B65717669AB8B1F7ED02022 ; reg IE4E0DDAB16DD8E970672626428251866 ; reg IE12D7FB0707DA0B72DA8BD64B6FAEFEB ;
reg I15C3BE43949B828A0A578329FE2EDE6B ; reg IE655D625D2EB067AC17967E600BE5FBD ; reg IABBE7E409672B3D3CE209351AE63C530 ;
reg I9962CDA8EE94C7BDFB23FE70815056E4 ; reg I7732946249B5963DFD9C95EC611A1D2C ; reg [6:0] I54D7451A32675B2129629BC41778D6D6 ;
reg [4:0] I8AC99AB880823B01C00D137F89AABEF8 ; reg [4:0] IF15E5692F18C2355720A228228564D0B ; reg IF8BC24CAD7E18C8A3A9A264889D5ECF8 ;
reg I9B8138DCE156F7C31EB5914EF01F183C ; reg [7:0] IB9A23596C80981B9B1CF7E12A76E71AC ; reg [4:0] I288715DFB3893A064D51571152559F12 ;
reg [2:0] I86B9557FA0123B8105E34300F4FCD447 ; reg [I63F1EFA9086319A16127622F3CE8B7D0 - 1:0] I3EC90F87E70407C2A46DA25A8CA9065B ;
reg [63:0] I9E40C3A9F9E3CDFC05F95566701DFB02 ; reg ICDFF33095CB0890DA2F167B63251EC67 ; reg IAE5BB83186BAD37A0D9A9B45FFE89934 ;
reg IB9889A1CC70F16308850E5AB5B9F99AF ; reg I5E1B26AB678FDA8FBEB1A0F43F21D9E4 ; reg [IDB9D60794264C5F8E5363941194A797B
- 1:0] I5B0AA124C4ADA63A064AF2CAFA1098FD ; reg [3:0] I93F6D99D18FD6FF40EF5AD5288D5C88E ; reg [63:0] I83F18730E4735495B20E29C862E672F1 ;
reg [13:0] I18D210808E8E4FD4E19269D50B767EF6 ; reg [10:0] I84B10D95B4B5E01F827E0D4D81BF476B ; reg [7:0] I539C1D01FC349447001EB93E17D37611 ;
reg [63:0] I2C5E6805594DFF3B9EB915045ABF7575 ; reg I41486045CC0DB09C489AD9C404A6348F ; reg [I63F1EFA9086319A16127622F3CE8B7D0
- 1:0] I909A2BB1C99AC88EE130F2C2B36CD5AB ; reg I893DF0D582AF0617B44879E65C202360 ; reg I2967174B668E2BB5A635A3F85DFF312B ;
reg I2212D954BC70C49C1F608E169DC873BC ; reg I5B3BB6CF473F793585E2668A9A7136C8 ; reg [ID7C7F9F2E39BEBEE2ACFA8040034E48D
- 1:0] IC7779D4175ADF3F75C21392F9E824B6D ; reg [1:0] IA6B00370F90E5BFE7B5D8852390CF107 ; reg [2:0] I369C3845EEBC3367BADAF446789A185D ;
reg I57E5F0C022683CA716D05ABE3408A469 ; reg IE7D8E2A0B7B7689804FFDF702BF724A6 ; reg I6F3C14B2AF4F4232F642DBEB36DCF09E ;
reg I33F9C80AA280FFCBE2A2CB54C2056CC5 ; reg [IDB9D60794264C5F8E5363941194A797B - 1:0] I5A4554E3FF0F3BAFC519CDF46237B987 ;
reg [31:0] I4A32ABD54816279F9EB5B44658C862FE ; reg [63:0] I074FD9C5AE408613B3750B75A6125486 ; reg I0EBD58BCF1D55F648B20B722C25EA4A8 ;
reg [10:0] I30D7DB78C2B62A00872F044F1A2F39A2 ; reg [10:0] IA934CBE3CC9AEBA0C32AA4C7EFA4954C ; reg [3:0] I13C229A5BDE90D9F920D8F4D218106DE ;
reg I037773E6A298229B4A19627ABA272E81 ; reg I36FECBB048E15937DC767259CBABEDCB ; wire [7:0] IC4C940842A3072C3A9C40616C6A213F2 ;
wire [4:0] IE8010EDEC4159FBD688A550900D0006D ; wire [2:0] I6345C4C803C15670FB2665AEA7AA4E33 ; wire IDEA2A0E5DD71C950358A21DDB6565B0A ;
wire I93FEA934E2F91A4D5E773376B9B26FED ; wire [63:0] IECBB27B02681BC7BD91D739A6D8B2975 ; wire [63:0] ID1BBB7750C0A323CA33FE43DEC09068C ;
wire IEDEC097EECBEE6B592219F6FEFFC7C2A ; wire I6FFEBECC6A03EE718A0503E2B1CA3AF0 ; wire [63:0] I1C0B5D2F7BB5720EB08D3892BAD2F2CA ;
 assign IC2E260CA356C994048CCB108C7E359D1 = IBFF7FD594C616C9EBAD12448149DA576 ; assign IE707B5D4A74BA1BD745B52E0C07932C0
= I5AF6C20F3950D58007B9C0BEA7C87198 ; assign I6E70C748D9C56227AB1182F36658AE5C = I0C9CC98CD774EDC9DF9AB513E5A8FB57 ;
assign I59B23598E8ADE1982F184EF67BEB0979 = I26F46DF735C89C3DA76F7F404A5F650F ; assign I33E409903692F5ECA2EC3553F9D1659E
= I533559C7D3A6FC7D4A2E49A02AFC9137 ; assign I437E57D42FB91B674CCBCC915BF9D653 = IF9A51F60DF053D68A5D57FECB5AB7ACB ;
assign I55AFDDE17B53D7F65849D39B02B07417 = I4A3B5CD6A0CBD18332DCF8ECB309CC92 ; assign I65FE2DB4E1CB5A488A45D60041AB5F64
= {I2931854F66F4E6D5E96ED7D73266F38E [7:0], I2931854F66F4E6D5E96ED7D73266F38E [15:8], I2931854F66F4E6D5E96ED7D73266F38E [23:16],
I2931854F66F4E6D5E96ED7D73266F38E [31:24]}; assign I0C796C206FE7060B578156D0110461EB = I83F18730E4735495B20E29C862E672F1 ;
assign IFC86A6522A8CA080A0DB7F384D9CE6FA = IE12D7FB0707DA0B72DA8BD64B6FAEFEB ; assign I484F77D7967D25736EB27A0ED76CCB5F
= I9C46AA186B65717669AB8B1F7ED02022 ; assign I7E0431D7F1A92C0ED1F030F36BF809B7 = IE4E0DDAB16DD8E970672626428251866 ;
assign I3E6965EC606FD6C2871F2C0993204C57 = I15C3BE43949B828A0A578329FE2EDE6B ; assign IFF25B820DFD457D71B32B130ABE5DA3F
= IE655D625D2EB067AC17967E600BE5FBD ; assign I20FA57C9A87CB2AA26088D9FA1743F70 = IABBE7E409672B3D3CE209351AE63C530 ;
assign I51C881E8B9B36D7A724BC7B8EC533957 = I511F58CE0ACA83EE959D1BF6C4EAFA7F ; assign ID3E7F4B58943229FEE6313A36B3F8693
= I7E9516402D6933186513EB5B37336278 ; assign I1FDEC1735547330C00A0B8DFE1FB10C3 = IA1EA4D4C05E159614ABC1E6D9CABE3BB ;
assign IBD6A65D48B4A68CA0D2A82F79053757B = I8916D921407646CE03BABA39B922EE09 ; assign I15EC78E3DE1101BFF2B227962683E113
= IEDEC097EECBEE6B592219F6FEFFC7C2A ; assign I7C4DADE2C05F6DCECCAF7AD6F7BF2FF8 = I2C5E6805594DFF3B9EB915045ABF7575 ;
assign IEEFA85D6664F09687B5CA591C701DC34 = I893DF0D582AF0617B44879E65C202360 ; assign ID4A284C76C6EABEEBA8E0AE18003FBAC
= I2212D954BC70C49C1F608E169DC873BC ; assign I6010C20131B976554A498745FEEEB580 = I5B3BB6CF473F793585E2668A9A7136C8 ;
assign I46E8CA15DC1E8B3B2200999A53029704 = IC7779D4175ADF3F75C21392F9E824B6D ; assign IEC45B60C7D1A49FFA84D3F5D121A2579
= IA6B00370F90E5BFE7B5D8852390CF107 ; assign I9AF46E2AA924FA7E0F5D7290324BABF9 = I369C3845EEBC3367BADAF446789A185D ;
assign I59D9A9A677978229C1F87AA1A3A0C304 = I57E5F0C022683CA716D05ABE3408A469 ; assign I9301CE4E9B877D08EDBD1584D6BE017A
= IE7D8E2A0B7B7689804FFDF702BF724A6 ; assign I51698892CBD372EE66AF3EA4D0ECE23F = I6F3C14B2AF4F4232F642DBEB36DCF09E ;
assign I1347408C9E757F34EA4D78F53447BD9B = I33F9C80AA280FFCBE2A2CB54C2056CC5 ; assign I2BE88607F3C31B47400F3A35E08B7EAD
= I5A4554E3FF0F3BAFC519CDF46237B987 ; assign I7D901091F9E0741061C75B54467D48A0 = I074FD9C5AE408613B3750B75A6125486 ;
assign I7AEBDB3D2CD4891A528BA81F5F54B20D = I0EBD58BCF1D55F648B20B722C25EA4A8 ; assign ID16819FEAA95700005E383E7DA0C8E13
= I30D7DB78C2B62A00872F044F1A2F39A2 ; assign IE0337CA803FBA20F38A0CD2A900C6534 = I11FD35FED78BCB8861FACB9A1E3A4C35 ;
assign I592A6A3BA99B09C24695C7A609F9053F = IC52F3B77F7E45A74323561D6A6F6028A ; assign I40EF39BB4F4F4A031C8FD1026EF53063
= I13C229A5BDE90D9F920D8F4D218106DE ; assign I42427E866FF31BC28E35C71EC172E26B = I037773E6A298229B4A19627ABA272E81 ;
assign I368749E68EAF9F462385FAD36180A9FE = I36FECBB048E15937DC767259CBABEDCB ;  assign IC4C940842A3072C3A9C40616C6A213F2
= (I511F58CE0ACA83EE959D1BF6C4EAFA7F & I9C46AA186B65717669AB8B1F7ED02022 ) ? I7E9516402D6933186513EB5B37336278 :
IFF5E23C5A17BB678C108274E28C56424 ; assign IE8010EDEC4159FBD688A550900D0006D = (I511F58CE0ACA83EE959D1BF6C4EAFA7F
& I9C46AA186B65717669AB8B1F7ED02022 ) ? IA1EA4D4C05E159614ABC1E6D9CABE3BB : IDE425A12275C43D9056DCF647A2D8258 ;
assign I6345C4C803C15670FB2665AEA7AA4E33 = (I511F58CE0ACA83EE959D1BF6C4EAFA7F & I9C46AA186B65717669AB8B1F7ED02022 )
? I8916D921407646CE03BABA39B922EE09 : I65B14714ECFCC218D3A788DF7696216B ; assign IDEA2A0E5DD71C950358A21DDB6565B0A
= (I7E600D684E83043922C1FE27CC6213E4 ) ? 1'b1 : 1'b0; assign IECBB27B02681BC7BD91D739A6D8B2975 = {I36824F33FF142FDE2AFE9BC4759DB690 [39:32],
I36824F33FF142FDE2AFE9BC4759DB690 [47:40], I36824F33FF142FDE2AFE9BC4759DB690 [55:48], I36824F33FF142FDE2AFE9BC4759DB690 [63:56],
I36824F33FF142FDE2AFE9BC4759DB690 [7:0], I36824F33FF142FDE2AFE9BC4759DB690 [15:8], I36824F33FF142FDE2AFE9BC4759DB690 [23:16],
I36824F33FF142FDE2AFE9BC4759DB690 [31:24]}; assign ID1BBB7750C0A323CA33FE43DEC09068C = {I9E40C3A9F9E3CDFC05F95566701DFB02 [39:32],
I9E40C3A9F9E3CDFC05F95566701DFB02 [47:40], I9E40C3A9F9E3CDFC05F95566701DFB02 [55:48], I9E40C3A9F9E3CDFC05F95566701DFB02 [63:56],
I9E40C3A9F9E3CDFC05F95566701DFB02 [7:0], I9E40C3A9F9E3CDFC05F95566701DFB02 [15:8], I9E40C3A9F9E3CDFC05F95566701DFB02 [23:16],
I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24]}; assign I93FEA934E2F91A4D5E773376B9B26FED = (I9C46AA186B65717669AB8B1F7ED02022
& IF5E7E4E58741BF3FE58442AB377ED57F ) | (IE12D7FB0707DA0B72DA8BD64B6FAEFEB & IFC18758E8987A9913FD94A5DFEE774E2 )
| (IE4E0DDAB16DD8E970672626428251866 & IF5B4924BEAEA6935367AC2739021882F ) | ((I15C3BE43949B828A0A578329FE2EDE6B
| IE655D625D2EB067AC17967E600BE5FBD ) & IDEA2A0E5DD71C950358A21DDB6565B0A ) | (IABBE7E409672B3D3CE209351AE63C530
& I7985A5A43CBBBC8E0D3FCFEE38DDF221 ); assign IEDEC097EECBEE6B592219F6FEFFC7C2A = IAE5BB83186BAD37A0D9A9B45FFE89934
| IB9889A1CC70F16308850E5AB5B9F99AF | I6FFEBECC6A03EE718A0503E2B1CA3AF0 | I5E1B26AB678FDA8FBEB1A0F43F21D9E4 ; assign
I6FFEBECC6A03EE718A0503E2B1CA3AF0 = (I84B10D95B4B5E01F827E0D4D81BF476B > 1) ? (I511F58CE0ACA83EE959D1BF6C4EAFA7F
& I07B0EBE8FBC21BDBE894D73C90EDC5AB ) : 1'b0; assign I1C0B5D2F7BB5720EB08D3892BAD2F2CA = {I3D6C771D05CA1A769E61302C086494B8 [7:0],
I3D6C771D05CA1A769E61302C086494B8 [15:8], I3D6C771D05CA1A769E61302C086494B8 [23:16], I3D6C771D05CA1A769E61302C086494B8 [31:24]};
 always @(*) begin IF15E5692F18C2355720A228228564D0B = I8AC99AB880823B01C00D137F89AABEF8 ; case (I8AC99AB880823B01C00D137F89AABEF8 )
I3662C12143A4A1B904AC8798CEEF0125 : begin if (I9F3623AEB414A15CECD2A8FD8791C79D > 1) IF15E5692F18C2355720A228228564D0B
= I257DF24B77C5CA85F676E7FFA065CE94 ; end I257DF24B77C5CA85F676E7FFA065CE94 : begin if (IA886199C0F7609B072DAE171DFC98CD8 )
IF15E5692F18C2355720A228228564D0B = I67E645B7D6135C108074CF368E9BB834 ; end I67E645B7D6135C108074CF368E9BB834 :
begin IF15E5692F18C2355720A228228564D0B = IFE893DBF9067A0DA39E179005AD783C4 ; end IFE893DBF9067A0DA39E179005AD783C4
: begin IF15E5692F18C2355720A228228564D0B = I56AC73D28E70D2F78200164359CC0E9A ; end I56AC73D28E70D2F78200164359CC0E9A
: begin if (IDA48F17DCE4BB1F6A04CBB23CCB4C3A5 == 0) IF15E5692F18C2355720A228228564D0B = I499DB4E92AEE1C97FE024F6FD8CDEB8A ;
end I499DB4E92AEE1C97FE024F6FD8CDEB8A : begin if (I93FEA934E2F91A4D5E773376B9B26FED ) if (I9962CDA8EE94C7BDFB23FE70815056E4 )
IF15E5692F18C2355720A228228564D0B = IC495D10CCC7452A18D769BDD99794652 ; else if (I511F58CE0ACA83EE959D1BF6C4EAFA7F )
IF15E5692F18C2355720A228228564D0B = IABEE3580E02F366EC5560A9CFC5CC953 ; else IF15E5692F18C2355720A228228564D0B =
I2D358EAE916810B434B6C76F7C7C5673 ; else IF15E5692F18C2355720A228228564D0B = IFAC7B411ECB5421590DDAA0B7B34F238 ;
end IABEE3580E02F366EC5560A9CFC5CC953 : begin if (ICDFF33095CB0890DA2F167B63251EC67 ) IF15E5692F18C2355720A228228564D0B
= I2D358EAE916810B434B6C76F7C7C5673 ; end I2D358EAE916810B434B6C76F7C7C5673 : begin IF15E5692F18C2355720A228228564D0B
= I174E152AA0198C30C57B401C947D37C1 ; end I174E152AA0198C30C57B401C947D37C1 : begin if (I511F58CE0ACA83EE959D1BF6C4EAFA7F )
begin if ((IA886199C0F7609B072DAE171DFC98CD8 == 1'b1) || ((IF4B2F356412545C21578876129150C2F == 1'b0) && (IA934CBE3CC9AEBA0C32AA4C7EFA4954C
== 1))) IF15E5692F18C2355720A228228564D0B = I29C10DD8DAC8AB31273614BA27A5E29C ; end else IF15E5692F18C2355720A228228564D0B
= I3C15F904BACDB851EFC4C548820E98B8 ; end I3C15F904BACDB851EFC4C548820E98B8 : begin if (I07B0EBE8FBC21BDBE894D73C90EDC5AB
& (IA934CBE3CC9AEBA0C32AA4C7EFA4954C == 1)) IF15E5692F18C2355720A228228564D0B = IF5A7A7CE92502E2DF9F0601605A38637 ;
end I29C10DD8DAC8AB31273614BA27A5E29C : begin if (I07B0EBE8FBC21BDBE894D73C90EDC5AB & (I84B10D95B4B5E01F827E0D4D81BF476B
== 0)) IF15E5692F18C2355720A228228564D0B = IF5A7A7CE92502E2DF9F0601605A38637 ; end IF5A7A7CE92502E2DF9F0601605A38637
: begin IF15E5692F18C2355720A228228564D0B = I5021A214EB457E909E76C621F6DD12B1 ; end I5021A214EB457E909E76C621F6DD12B1
: begin if (I7FA4C54BD6B551C794EE0EA588CBD4C7 ) IF15E5692F18C2355720A228228564D0B = I05E305FFF5B6CDE122F8935EE521D523 ;
else IF15E5692F18C2355720A228228564D0B = I3662C12143A4A1B904AC8798CEEF0125 ; end I05E305FFF5B6CDE122F8935EE521D523
: begin if (I9F4F7E2C4A4A8FB2780021EDF6E4ADEF ) IF15E5692F18C2355720A228228564D0B = I3662C12143A4A1B904AC8798CEEF0125 ;
end IFAC7B411ECB5421590DDAA0B7B34F238 : begin if (I511F58CE0ACA83EE959D1BF6C4EAFA7F ) begin if (ICDFF33095CB0890DA2F167B63251EC67 )
IF15E5692F18C2355720A228228564D0B = I248DCDE6260EE21AB43E9E1EF6D603EF ; end else begin if (I9962CDA8EE94C7BDFB23FE70815056E4 )
IF15E5692F18C2355720A228228564D0B = I6EA1237B063AFA6C82E354D0001BEF41 ; else IF15E5692F18C2355720A228228564D0B =
IF5A7A7CE92502E2DF9F0601605A38637 ; end end I248DCDE6260EE21AB43E9E1EF6D603EF : begin if ((IEDEC097EECBEE6B592219F6FEFFC7C2A )
&& (I84B10D95B4B5E01F827E0D4D81BF476B == 1)) if (I9962CDA8EE94C7BDFB23FE70815056E4 ) IF15E5692F18C2355720A228228564D0B
= I6EA1237B063AFA6C82E354D0001BEF41 ; else IF15E5692F18C2355720A228228564D0B = IF5A7A7CE92502E2DF9F0601605A38637 ;
end IC495D10CCC7452A18D769BDD99794652 : begin if (ICB518A59CAE27DDB6398AB22F5D74259 > 2) IF15E5692F18C2355720A228228564D0B
= I6EA1237B063AFA6C82E354D0001BEF41 ; end IEAE55E29AC7D8EC5093BF4C91D5CFFCE : begin if (I2967174B668E2BB5A635A3F85DFF312B )
IF15E5692F18C2355720A228228564D0B = I2D358EAE916810B434B6C76F7C7C5673 ; end I6EA1237B063AFA6C82E354D0001BEF41 :
begin IF15E5692F18C2355720A228228564D0B = I070181DB2ED3EDD3633DB4E93B8E42A5 ; end I070181DB2ED3EDD3633DB4E93B8E42A5
: begin IF15E5692F18C2355720A228228564D0B = I2263EE3B1CDD9957F685B729A9639643 ; end I2263EE3B1CDD9957F685B729A9639643
: begin if (I7732946249B5963DFD9C95EC611A1D2C ) IF15E5692F18C2355720A228228564D0B = IF5A7A7CE92502E2DF9F0601605A38637 ;
else if (I511F58CE0ACA83EE959D1BF6C4EAFA7F ) IF15E5692F18C2355720A228228564D0B = IABEE3580E02F366EC5560A9CFC5CC953 ;
else IF15E5692F18C2355720A228228564D0B = IEAE55E29AC7D8EC5093BF4C91D5CFFCE ; end default : begin end endcase end
 always @(posedge ICCFB0F435B37370076102F325BC08D20 or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin : I50905559064282CED274D62360FCE175
if (~I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin I11FD35FED78BCB8861FACB9A1E3A4C35 <= 4'hf; IC52F3B77F7E45A74323561D6A6F6028A
<= 4'hf; I0FF03F7D70F3047C91A55F9744DDD7AE <= 1'b0; IAC85A6B0EE1F3079B60C115CB476DF06 <= 12'b0; I71DBDE411F9CED520FD43A4EF5CBD656
<= 9'b0; IBFF7FD594C616C9EBAD12448149DA576 <= 8'b0; I0C9CC98CD774EDC9DF9AB513E5A8FB57 <= 1'b0; I26F46DF735C89C3DA76F7F404A5F650F
<= 1'b0; I5AF6C20F3950D58007B9C0BEA7C87198 <= 8'b0; I533559C7D3A6FC7D4A2E49A02AFC9137 <= 1'b0; IF9A51F60DF053D68A5D57FECB5AB7ACB
<= 1'b0; I916551CA30E7A94681BA2B3415BF85FA <= 1'b0; I4A3B5CD6A0CBD18332DCF8ECB309CC92 <= 1'b0; I2931854F66F4E6D5E96ED7D73266F38E
<= 64'b0; IDA48F17DCE4BB1F6A04CBB23CCB4C3A5 <= {I15DA3B10E1E0658D2D01B744DF560903 {1'b0}}; IC93C4C87277AF77C73E35A77E14FC4B1
<= 1'b0; I54BE80AB8C90F3E5819921EF5354732A <= 1'b0; I7FA4C54BD6B551C794EE0EA588CBD4C7 <= 1'b0; I511F58CE0ACA83EE959D1BF6C4EAFA7F
<= 1'b0; IF4B2F356412545C21578876129150C2F <= 1'b0; I7E9516402D6933186513EB5B37336278 <= 8'b0; IA1EA4D4C05E159614ABC1E6D9CABE3BB
<= 5'b0; I8916D921407646CE03BABA39B922EE09 <= 3'b0; I9C46AA186B65717669AB8B1F7ED02022 <= 1'b0; IE4E0DDAB16DD8E970672626428251866
<= 1'b0; IE12D7FB0707DA0B72DA8BD64B6FAEFEB <= 1'b0; I15C3BE43949B828A0A578329FE2EDE6B <= 1'b0; IE655D625D2EB067AC17967E600BE5FBD
<= 1'b0; IABBE7E409672B3D3CE209351AE63C530 <= 1'b0; I9962CDA8EE94C7BDFB23FE70815056E4 <= 1'b0; I7732946249B5963DFD9C95EC611A1D2C
<= 1'b0; I54D7451A32675B2129629BC41778D6D6 <= 7'b0; I8AC99AB880823B01C00D137F89AABEF8 <= I3662C12143A4A1B904AC8798CEEF0125 ;
IF8BC24CAD7E18C8A3A9A264889D5ECF8 <= 1'b0; I9B8138DCE156F7C31EB5914EF01F183C <= 1'b0; IB9A23596C80981B9B1CF7E12A76E71AC
<= 8'b0; I288715DFB3893A064D51571152559F12 <= 5'b0; I86B9557FA0123B8105E34300F4FCD447 <= 3'b0; I3EC90F87E70407C2A46DA25A8CA9065B
<= {I63F1EFA9086319A16127622F3CE8B7D0 {1'b0}}; I9E40C3A9F9E3CDFC05F95566701DFB02 <= 64'b0; ICDFF33095CB0890DA2F167B63251EC67
<= 1'b0; IAE5BB83186BAD37A0D9A9B45FFE89934 <= 1'b0; IB9889A1CC70F16308850E5AB5B9F99AF <= 1'b0; I5E1B26AB678FDA8FBEB1A0F43F21D9E4
<= 1'b0; I5B0AA124C4ADA63A064AF2CAFA1098FD <= {IDB9D60794264C5F8E5363941194A797B {1'b0}}; I93F6D99D18FD6FF40EF5AD5288D5C88E
<= 4'b0; I83F18730E4735495B20E29C862E672F1 <= 64'b0; I18D210808E8E4FD4E19269D50B767EF6 <= 14'b0; I84B10D95B4B5E01F827E0D4D81BF476B
<= 11'b0; I539C1D01FC349447001EB93E17D37611 <= 8'b0; I5B3BB6CF473F793585E2668A9A7136C8 <= 1'b0; I2C5E6805594DFF3B9EB915045ABF7575
<= 64'b0; I41486045CC0DB09C489AD9C404A6348F <= 1'b0; I909A2BB1C99AC88EE130F2C2B36CD5AB <= {I63F1EFA9086319A16127622F3CE8B7D0 {1'b0}};
I893DF0D582AF0617B44879E65C202360 <= 1'b0; I2967174B668E2BB5A635A3F85DFF312B <= 1'b0; I2212D954BC70C49C1F608E169DC873BC
<= 1'b0; IC7779D4175ADF3F75C21392F9E824B6D <= {ID7C7F9F2E39BEBEE2ACFA8040034E48D {1'b0}}; IA6B00370F90E5BFE7B5D8852390CF107
<= 2'b0; I369C3845EEBC3367BADAF446789A185D <= 3'b0; I57E5F0C022683CA716D05ABE3408A469 <= 1'b0; IE7D8E2A0B7B7689804FFDF702BF724A6
<= 1'b0; I6F3C14B2AF4F4232F642DBEB36DCF09E <= 1'b0; I33F9C80AA280FFCBE2A2CB54C2056CC5 <= 1'b0; I5A4554E3FF0F3BAFC519CDF46237B987
<= {IDB9D60794264C5F8E5363941194A797B {1'b0}}; I4A32ABD54816279F9EB5B44658C862FE <= {32{1'b0}}; I074FD9C5AE408613B3750B75A6125486
<= 64'b0; IA934CBE3CC9AEBA0C32AA4C7EFA4954C <= 12'b0; I13C229A5BDE90D9F920D8F4D218106DE <= 4'b0; I037773E6A298229B4A19627ABA272E81
<= 1'b0; I0EBD58BCF1D55F648B20B722C25EA4A8 <= 1'b0; I30D7DB78C2B62A00872F044F1A2F39A2 <= {11{1'b0}}; I36FECBB048E15937DC767259CBABEDCB
<= 1'b0; end else begin I4A3B5CD6A0CBD18332DCF8ECB309CC92 <= IA886199C0F7609B072DAE171DFC98CD8 & I916551CA30E7A94681BA2B3415BF85FA ;
I2931854F66F4E6D5E96ED7D73266F38E <= I36824F33FF142FDE2AFE9BC4759DB690 ; I54BE80AB8C90F3E5819921EF5354732A <= I93AE636CE82DE94CB11ACCF59F8C2254 ;
I8AC99AB880823B01C00D137F89AABEF8 <= IF15E5692F18C2355720A228228564D0B ; I3EC90F87E70407C2A46DA25A8CA9065B <= I9F3623AEB414A15CECD2A8FD8791C79D ;
ICDFF33095CB0890DA2F167B63251EC67 <= 1'b1;  IAE5BB83186BAD37A0D9A9B45FFE89934 <= 1'b0; IB9889A1CC70F16308850E5AB5B9F99AF
<= 1'b0; I5E1B26AB678FDA8FBEB1A0F43F21D9E4 <= 1'b0; I909A2BB1C99AC88EE130F2C2B36CD5AB <= ICB518A59CAE27DDB6398AB22F5D74259 ;
I893DF0D582AF0617B44879E65C202360 <= 1'b0; I2967174B668E2BB5A635A3F85DFF312B <= (I909A2BB1C99AC88EE130F2C2B36CD5AB
>= IA934CBE3CC9AEBA0C32AA4C7EFA4954C ) ? 1'b1 : 1'b0; I2212D954BC70C49C1F608E169DC873BC <= 1'b0; I0EBD58BCF1D55F648B20B722C25EA4A8
<= 1'b0; if (IA886199C0F7609B072DAE171DFC98CD8 == 1'b1) I9E40C3A9F9E3CDFC05F95566701DFB02 <= I36824F33FF142FDE2AFE9BC4759DB690 ;
case (I8AC99AB880823B01C00D137F89AABEF8 ) I3662C12143A4A1B904AC8798CEEF0125 : begin I916551CA30E7A94681BA2B3415BF85FA
<= 1'b0; IB9889A1CC70F16308850E5AB5B9F99AF <= (I9F3623AEB414A15CECD2A8FD8791C79D > 1) ? 1'b1 : 1'b0; end I257DF24B77C5CA85F676E7FFA065CE94
: begin IDA48F17DCE4BB1F6A04CBB23CCB4C3A5 <= I15DA3B10E1E0658D2D01B744DF560903 - 1; I9E40C3A9F9E3CDFC05F95566701DFB02
<= I36824F33FF142FDE2AFE9BC4759DB690 ; IB9889A1CC70F16308850E5AB5B9F99AF <= 1'b1; I83F18730E4735495B20E29C862E672F1
<= {64{1'b0}}; I893DF0D582AF0617B44879E65C202360 <= 1'b0; end I67E645B7D6135C108074CF368E9BB834 : begin I11FD35FED78BCB8861FACB9A1E3A4C35
<= I9E40C3A9F9E3CDFC05F95566701DFB02 [35:32]; IC52F3B77F7E45A74323561D6A6F6028A <= I9E40C3A9F9E3CDFC05F95566701DFB02 [39:36];
I7FA4C54BD6B551C794EE0EA588CBD4C7 <= 1'b0; I511F58CE0ACA83EE959D1BF6C4EAFA7F <= I9E40C3A9F9E3CDFC05F95566701DFB02 [30];
IF4B2F356412545C21578876129150C2F <= I9E40C3A9F9E3CDFC05F95566701DFB02 [29]; IB9A23596C80981B9B1CF7E12A76E71AC <=
I9E40C3A9F9E3CDFC05F95566701DFB02 [63:56]; I288715DFB3893A064D51571152559F12 <= I9E40C3A9F9E3CDFC05F95566701DFB02 [55:51];
I86B9557FA0123B8105E34300F4FCD447 <= I9E40C3A9F9E3CDFC05F95566701DFB02 [50:48]; I18D210808E8E4FD4E19269D50B767EF6
<= I9E40C3A9F9E3CDFC05F95566701DFB02 [23:10]; I84B10D95B4B5E01F827E0D4D81BF476B <= {1'b0, I9E40C3A9F9E3CDFC05F95566701DFB02 [10:0]};
I84B10D95B4B5E01F827E0D4D81BF476B <= {((I9E40C3A9F9E3CDFC05F95566701DFB02 [9:0] == 0) ? 1'b1 : 1'b0), I9E40C3A9F9E3CDFC05F95566701DFB02 [9:0]};
I539C1D01FC349447001EB93E17D37611 <= I9E40C3A9F9E3CDFC05F95566701DFB02 [47:40]; I9C46AA186B65717669AB8B1F7ED02022
<= ((I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I81D26620360085DCC2783D5734873451 ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24]
== IA3187A41E33086C9DA805D8C67004992 )) ? 1'b1 : 1'b0; IE4E0DDAB16DD8E970672626428251866 <= ((I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24]
== I2C8281C2456BAC869C04372CE6A7C50E ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I8CD6057CFBD7215340EF60C41A0C63EC ))
? 1'b1 : 1'b0; IE12D7FB0707DA0B72DA8BD64B6FAEFEB <= ((I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I6A62FD6104E281B8714322DB8CCB5FE3 )
|| (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I85B0192F2AC4464C88E2C93352FE6696 ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24]
== I78DDE5821936F928E302A8BA3C3138EE ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I41F249A62806D544C38454CA2D10750D ))
? 1'b1 : 1'b0; I15C3BE43949B828A0A578329FE2EDE6B <= ((I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I34EF8B0D0058C1876C19361DBBAC62DC )
|| (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == IB83A8F7EA6693A633C486F9CA18003BB )) ? 1'b1 : 1'b0; IE655D625D2EB067AC17967E600BE5FBD
<= ((I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I8F0EB88EC813DC0B3105F31BABD34B79 ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24]
== I877B2A234FC10EC8A4A2F0A90F6EAE6C ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == IEC10F95DD42CAF869EFB03BDF59BE8EB )
|| (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I2E664E814B6AA2CBCE57FBCE2A354435 )) ? 1'b1 : 1'b0; IABBE7E409672B3D3CE209351AE63C530
<= (((I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] & 8'hf0) == IBC983AF54FD90EA2AA9E3DD139A3B818 ) || ((I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24]
& 8'hf0) == I361F321AEF89DD0EF2CEAC65B8B042D8 )) ? 1'b1 : 1'b0; I9962CDA8EE94C7BDFB23FE70815056E4 <= ((I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24]
== I8F0EB88EC813DC0B3105F31BABD34B79 ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I877B2A234FC10EC8A4A2F0A90F6EAE6C )
|| (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I81D26620360085DCC2783D5734873451 ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24]
== IA3187A41E33086C9DA805D8C67004992 ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I2C8281C2456BAC869C04372CE6A7C50E )
|| (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == I8CD6057CFBD7215340EF60C41A0C63EC ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24]
== I34EF8B0D0058C1876C19361DBBAC62DC ) || (I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24] == IB83A8F7EA6693A633C486F9CA18003BB ))
? 1'b1 : 1'b0; end IFE893DBF9067A0DA39E179005AD783C4 : begin IC52F3B77F7E45A74323561D6A6F6028A <= (I84B10D95B4B5E01F827E0D4D81BF476B
< 2) ? {4{1'b0}} : IC52F3B77F7E45A74323561D6A6F6028A ; I71DBDE411F9CED520FD43A4EF5CBD656 <= (I84B10D95B4B5E01F827E0D4D81BF476B [1:0]
== 2'b00) ? I84B10D95B4B5E01F827E0D4D81BF476B [10:2] : I84B10D95B4B5E01F827E0D4D81BF476B [10:2] + 1; I7E9516402D6933186513EB5B37336278
<= I9E40C3A9F9E3CDFC05F95566701DFB02 [31:24]; IA1EA4D4C05E159614ABC1E6D9CABE3BB <= I9E40C3A9F9E3CDFC05F95566701DFB02 [23:19];
I8916D921407646CE03BABA39B922EE09 <= I9E40C3A9F9E3CDFC05F95566701DFB02 [18:16]; IF8BC24CAD7E18C8A3A9A264889D5ECF8
<= (I15C3BE43949B828A0A578329FE2EDE6B | I9C46AA186B65717669AB8B1F7ED02022 | IE4E0DDAB16DD8E970672626428251866 )
? 1'b0 : ((I84B10D95B4B5E01F827E0D4D81BF476B > 1) ? ((~IF4B2F356412545C21578876129150C2F & ~I83F18730E4735495B20E29C862E672F1 [2])
| (IF4B2F356412545C21578876129150C2F & I83F18730E4735495B20E29C862E672F1 [2])) : 1'b0); IC7779D4175ADF3F75C21392F9E824B6D
<= {ID7C7F9F2E39BEBEE2ACFA8040034E48D {1'b0}}; I30D7DB78C2B62A00872F044F1A2F39A2 <= I84B10D95B4B5E01F827E0D4D81BF476B ;
IA934CBE3CC9AEBA0C32AA4C7EFA4954C <= I84B10D95B4B5E01F827E0D4D81BF476B ; if (I9C46AA186B65717669AB8B1F7ED02022 |
IE4E0DDAB16DD8E970672626428251866 ) begin I83F18730E4735495B20E29C862E672F1 [31:0] <= {17'b0, I9E40C3A9F9E3CDFC05F95566701DFB02 [18:16],
I9E40C3A9F9E3CDFC05F95566701DFB02 [11:0]}; I83F18730E4735495B20E29C862E672F1 [63:32] <= {32{1'b0}}; end else begin
I83F18730E4735495B20E29C862E672F1 <= (IF4B2F356412545C21578876129150C2F ) ? I9E40C3A9F9E3CDFC05F95566701DFB02 :
{{32{1'b0}}, I9E40C3A9F9E3CDFC05F95566701DFB02 [31:0]}; end case (IC52F3B77F7E45A74323561D6A6F6028A ) 4'b0100, 4'b0101,
4'b0110, 4'b0111 : case (I11FD35FED78BCB8861FACB9A1E3A4C35 ) 4'b0010, 4'b0110, 4'b1010, 4'b1110 : I93F6D99D18FD6FF40EF5AD5288D5C88E
<= 4'd2; 4'b0100, 4'b1100 : I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd3; 4'b1000 : I93F6D99D18FD6FF40EF5AD5288D5C88E
<= 4'd4; default I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd1; endcase 4'b0010, 4'b0011 : case (I11FD35FED78BCB8861FACB9A1E3A4C35 )
4'b0010, 4'b0110, 4'b1010, 4'b1110 : I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd3; 4'b0100, 4'b1100 : I93F6D99D18FD6FF40EF5AD5288D5C88E
<= 4'd4; 4'b1000 : I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd5; default I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd2;
endcase 4'b0001 : case (I11FD35FED78BCB8861FACB9A1E3A4C35 ) 4'b0010, 4'b0110, 4'b1010, 4'b1110 : I93F6D99D18FD6FF40EF5AD5288D5C88E
<= 4'd4; 4'b0100, 4'b1100 : I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd5; 4'b1000 : I93F6D99D18FD6FF40EF5AD5288D5C88E
<= 4'd6; default I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd3; endcase 4'b0000 : case (I11FD35FED78BCB8861FACB9A1E3A4C35 )
4'b0000, 4'b0001, 4'b0010, 4'b0100, 4'b1000 : I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd3; 4'b0011, 4'b0110, 4'b1100
: I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd2; 4'b0101, 4'b0111, 4'b1010, 4'b1110 : I93F6D99D18FD6FF40EF5AD5288D5C88E
<= 4'd1; default I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd0; endcase default case (I11FD35FED78BCB8861FACB9A1E3A4C35 )
4'b0010, 4'b0110, 4'b1010, 4'b1110 : I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd1; 4'b0100, 4'b1100 : I93F6D99D18FD6FF40EF5AD5288D5C88E
<= 4'd2; 4'b1000 : I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd3; default I93F6D99D18FD6FF40EF5AD5288D5C88E <= 4'd0;
endcase endcase end I56AC73D28E70D2F78200164359CC0E9A : begin I0FF03F7D70F3047C91A55F9744DDD7AE <= (IB9A23596C80981B9B1CF7E12A76E71AC
== IFF5E23C5A17BB678C108274E28C56424 ) ? 1'b1 : 1'b0; IC93C4C87277AF77C73E35A77E14FC4B1 <= (I288715DFB3893A064D51571152559F12
== IDE425A12275C43D9056DCF647A2D8258 ) ? 1'b1 : 1'b0; if (IDA48F17DCE4BB1F6A04CBB23CCB4C3A5 ) IDA48F17DCE4BB1F6A04CBB23CCB4C3A5
<= IDA48F17DCE4BB1F6A04CBB23CCB4C3A5 - 1; end I499DB4E92AEE1C97FE024F6FD8CDEB8A : begin IAC85A6B0EE1F3079B60C115CB476DF06
<= {I30D7DB78C2B62A00872F044F1A2F39A2 [9:0], 2'b00} - I93F6D99D18FD6FF40EF5AD5288D5C88E ; I916551CA30E7A94681BA2B3415BF85FA
<= IE12D7FB0707DA0B72DA8BD64B6FAEFEB & ((I7E9516402D6933186513EB5B37336278 == IFF5E23C5A17BB678C108274E28C56424 )
? 1'b1 : 1'b0) & ((IA1EA4D4C05E159614ABC1E6D9CABE3BB == IDE425A12275C43D9056DCF647A2D8258 ) ? 1'b1 : 1'b0); I7732946249B5963DFD9C95EC611A1D2C
<= ~I93FEA934E2F91A4D5E773376B9B26FED ; I5B0AA124C4ADA63A064AF2CAFA1098FD <= (IE655D625D2EB067AC17967E600BE5FBD
| I15C3BE43949B828A0A578329FE2EDE6B ) ? I7E600D684E83043922C1FE27CC6213E4 : {IDB9D60794264C5F8E5363941194A797B {1'b0}};
end I2D358EAE916810B434B6C76F7C7C5673 : begin IAE5BB83186BAD37A0D9A9B45FFE89934 <= ((I84B10D95B4B5E01F827E0D4D81BF476B
> 1) || IF4B2F356412545C21578876129150C2F ) ? I511F58CE0ACA83EE959D1BF6C4EAFA7F : 1'b0; end I174E152AA0198C30C57B401C947D37C1 :
begin if ((IA886199C0F7609B072DAE171DFC98CD8 == 1'b1) || (I511F58CE0ACA83EE959D1BF6C4EAFA7F == 1'b0) || ((IF4B2F356412545C21578876129150C2F
== 1'b0) && (IA934CBE3CC9AEBA0C32AA4C7EFA4954C == 1))) begin IA6B00370F90E5BFE7B5D8852390CF107 <= I6768A159F7F57847F9535CB8B8B382D8 ;
I57E5F0C022683CA716D05ABE3408A469 <= I9C46AA186B65717669AB8B1F7ED02022 ; IE7D8E2A0B7B7689804FFDF702BF724A6 <= IE4E0DDAB16DD8E970672626428251866 ;
I6F3C14B2AF4F4232F642DBEB36DCF09E <= IE12D7FB0707DA0B72DA8BD64B6FAEFEB ; I369C3845EEBC3367BADAF446789A185D <= (I84B10D95B4B5E01F827E0D4D81BF476B
== 1) ? IEE94C2462F89091D3C62992327532D1E : (((I84B10D95B4B5E01F827E0D4D81BF476B == 2) && IF4B2F356412545C21578876129150C2F )
? IEE94C2462F89091D3C62992327532D1E : I88A97019335E3F57955B11E67DFFCD65 ); I33F9C80AA280FFCBE2A2CB54C2056CC5 <=
IABBE7E409672B3D3CE209351AE63C530 ; I5A4554E3FF0F3BAFC519CDF46237B987 <= I5B0AA124C4ADA63A064AF2CAFA1098FD ; I037773E6A298229B4A19627ABA272E81
<= 1'b1; I0EBD58BCF1D55F648B20B722C25EA4A8 <= 1'b1; I36FECBB048E15937DC767259CBABEDCB <= I511F58CE0ACA83EE959D1BF6C4EAFA7F ;
if (IE12D7FB0707DA0B72DA8BD64B6FAEFEB ) IC7779D4175ADF3F75C21392F9E824B6D [14:0] <= {I86B9557FA0123B8105E34300F4FCD447 ,
I83F18730E4735495B20E29C862E672F1 [11:2], 2'b00}; else IC7779D4175ADF3F75C21392F9E824B6D <= {I83F18730E4735495B20E29C862E672F1 [ID7C7F9F2E39BEBEE2ACFA8040034E48D
- 1:2], 2'b00}; if (I511F58CE0ACA83EE959D1BF6C4EAFA7F ) begin if (I9C46AA186B65717669AB8B1F7ED02022 | IE4E0DDAB16DD8E970672626428251866 )
I074FD9C5AE408613B3750B75A6125486 <= {{32{1'b0}}, ID1BBB7750C0A323CA33FE43DEC09068C [63:32]}; else if (I15C3BE43949B828A0A578329FE2EDE6B )
I074FD9C5AE408613B3750B75A6125486 <= {ID1BBB7750C0A323CA33FE43DEC09068C [63:32], ID1BBB7750C0A323CA33FE43DEC09068C [31:0]};
else if (IF4B2F356412545C21578876129150C2F ) I074FD9C5AE408613B3750B75A6125486 <= (I83F18730E4735495B20E29C862E672F1 [2])
? {IECBB27B02681BC7BD91D739A6D8B2975 [31:0], {32{1'b0}}} : IECBB27B02681BC7BD91D739A6D8B2975 ; else I074FD9C5AE408613B3750B75A6125486
<= (I83F18730E4735495B20E29C862E672F1 [2]) ? {ID1BBB7750C0A323CA33FE43DEC09068C [63:32], {32{1'b0}}} : {IECBB27B02681BC7BD91D739A6D8B2975 [31:0],
ID1BBB7750C0A323CA33FE43DEC09068C [63:32]}; end if (I9C46AA186B65717669AB8B1F7ED02022 | IE4E0DDAB16DD8E970672626428251866 )
begin I84B10D95B4B5E01F827E0D4D81BF476B <= I84B10D95B4B5E01F827E0D4D81BF476B - 1; I13C229A5BDE90D9F920D8F4D218106DE
<= {{4{1'b0}}, I11FD35FED78BCB8861FACB9A1E3A4C35 }; end else if (I15C3BE43949B828A0A578329FE2EDE6B ) begin I84B10D95B4B5E01F827E0D4D81BF476B
<= I84B10D95B4B5E01F827E0D4D81BF476B - 1; I13C229A5BDE90D9F920D8F4D218106DE <= (I83F18730E4735495B20E29C862E672F1 [2])
? {I11FD35FED78BCB8861FACB9A1E3A4C35 , {4{1'b0}}} : {{4{1'b0}}, I11FD35FED78BCB8861FACB9A1E3A4C35 }; end else begin
I84B10D95B4B5E01F827E0D4D81BF476B <= (I83F18730E4735495B20E29C862E672F1 [2]) ? I84B10D95B4B5E01F827E0D4D81BF476B
- 1 : ((I84B10D95B4B5E01F827E0D4D81BF476B > 1) ? I84B10D95B4B5E01F827E0D4D81BF476B - 2 : I84B10D95B4B5E01F827E0D4D81BF476B
- 1); I13C229A5BDE90D9F920D8F4D218106DE <= (I83F18730E4735495B20E29C862E672F1 [2]) ? {I11FD35FED78BCB8861FACB9A1E3A4C35 ,
{4{1'b0}}} : ((I84B10D95B4B5E01F827E0D4D81BF476B > 2) ? {{4{1'b1}}, I11FD35FED78BCB8861FACB9A1E3A4C35 } : {IC52F3B77F7E45A74323561D6A6F6028A ,
I11FD35FED78BCB8861FACB9A1E3A4C35 }); end end end I3C15F904BACDB851EFC4C548820E98B8 : begin I2212D954BC70C49C1F608E169DC873BC
<= I07B0EBE8FBC21BDBE894D73C90EDC5AB ; if (I07B0EBE8FBC21BDBE894D73C90EDC5AB ) begin I41486045CC0DB09C489AD9C404A6348F
<= 1'b0; I893DF0D582AF0617B44879E65C202360 <= (I369C3845EEBC3367BADAF446789A185D == IEE94C2462F89091D3C62992327532D1E )
? 1'b1 : 1'b0; I369C3845EEBC3367BADAF446789A185D <= (IA934CBE3CC9AEBA0C32AA4C7EFA4954C == 2) ? IEE94C2462F89091D3C62992327532D1E
: I88A97019335E3F57955B11E67DFFCD65 ; I4A32ABD54816279F9EB5B44658C862FE <= I1C0B5D2F7BB5720EB08D3892BAD2F2CA [63:32];
I13C229A5BDE90D9F920D8F4D218106DE <= 4'b1111; IA934CBE3CC9AEBA0C32AA4C7EFA4954C <= (I41486045CC0DB09C489AD9C404A6348F )
? IA934CBE3CC9AEBA0C32AA4C7EFA4954C - 1 : ((IA934CBE3CC9AEBA0C32AA4C7EFA4954C > 1) ? IA934CBE3CC9AEBA0C32AA4C7EFA4954C
- 2 : IA934CBE3CC9AEBA0C32AA4C7EFA4954C - 1); if (I9B8138DCE156F7C31EB5914EF01F183C ) if (I9C46AA186B65717669AB8B1F7ED02022
| IE4E0DDAB16DD8E970672626428251866 ) I2C5E6805594DFF3B9EB915045ABF7575 <= {I2C5E6805594DFF3B9EB915045ABF7575 [63:32],
I1C0B5D2F7BB5720EB08D3892BAD2F2CA [31:0]}; else if (I15C3BE43949B828A0A578329FE2EDE6B ) I2C5E6805594DFF3B9EB915045ABF7575
<= {((I54D7451A32675B2129629BC41778D6D6 [2]) ? I1C0B5D2F7BB5720EB08D3892BAD2F2CA [63:32] : I1C0B5D2F7BB5720EB08D3892BAD2F2CA [31:0]),
I2C5E6805594DFF3B9EB915045ABF7575 [31:0]}; else if (I41486045CC0DB09C489AD9C404A6348F ) I2C5E6805594DFF3B9EB915045ABF7575
<= {((I54D7451A32675B2129629BC41778D6D6 [2]) ? I1C0B5D2F7BB5720EB08D3892BAD2F2CA [63:32] : I1C0B5D2F7BB5720EB08D3892BAD2F2CA [31:0]),
I2C5E6805594DFF3B9EB915045ABF7575 [31:0]}; else I2C5E6805594DFF3B9EB915045ABF7575 <= (IF8BC24CAD7E18C8A3A9A264889D5ECF8 )
? {I1C0B5D2F7BB5720EB08D3892BAD2F2CA [31:0], I2C5E6805594DFF3B9EB915045ABF7575 [31:0]} : I1C0B5D2F7BB5720EB08D3892BAD2F2CA ;
else I2C5E6805594DFF3B9EB915045ABF7575 <= {64{1'b1}}; if (I369C3845EEBC3367BADAF446789A185D == IEE94C2462F89091D3C62992327532D1E )
begin IC7779D4175ADF3F75C21392F9E824B6D <= {ID7C7F9F2E39BEBEE2ACFA8040034E48D {1'b0}}; I074FD9C5AE408613B3750B75A6125486
<= 64'b0; IA6B00370F90E5BFE7B5D8852390CF107 <= 2'b0; I369C3845EEBC3367BADAF446789A185D <= 3'b0; I57E5F0C022683CA716D05ABE3408A469
<= 1'b0; IE7D8E2A0B7B7689804FFDF702BF724A6 <= 1'b0; I6F3C14B2AF4F4232F642DBEB36DCF09E <= 1'b0; I33F9C80AA280FFCBE2A2CB54C2056CC5
<= 1'b0; I5A4554E3FF0F3BAFC519CDF46237B987 <= {IDB9D60794264C5F8E5363941194A797B {1'b0}}; I13C229A5BDE90D9F920D8F4D218106DE
<= 4'b0; I037773E6A298229B4A19627ABA272E81 <= 1'b0; I36FECBB048E15937DC767259CBABEDCB <= 1'b0; end end end I29C10DD8DAC8AB31273614BA27A5E29C
: begin if (IEDEC097EECBEE6B592219F6FEFFC7C2A ) I9E40C3A9F9E3CDFC05F95566701DFB02 <= I36824F33FF142FDE2AFE9BC4759DB690 ;
if (I07B0EBE8FBC21BDBE894D73C90EDC5AB ) begin I84B10D95B4B5E01F827E0D4D81BF476B <= (I84B10D95B4B5E01F827E0D4D81BF476B
> 1) ? I84B10D95B4B5E01F827E0D4D81BF476B - 2 : I84B10D95B4B5E01F827E0D4D81BF476B - 1; if (I369C3845EEBC3367BADAF446789A185D
== IEE94C2462F89091D3C62992327532D1E ) begin IC7779D4175ADF3F75C21392F9E824B6D <= {ID7C7F9F2E39BEBEE2ACFA8040034E48D {1'b0}};
I074FD9C5AE408613B3750B75A6125486 <= {64{1'b0}}; IA6B00370F90E5BFE7B5D8852390CF107 <= 2'b0; I369C3845EEBC3367BADAF446789A185D
<= 3'b0; I57E5F0C022683CA716D05ABE3408A469 <= 1'b0; IE7D8E2A0B7B7689804FFDF702BF724A6 <= 1'b0; I6F3C14B2AF4F4232F642DBEB36DCF09E
<= 1'b0; I33F9C80AA280FFCBE2A2CB54C2056CC5 <= 1'b0; I5A4554E3FF0F3BAFC519CDF46237B987 <= {IDB9D60794264C5F8E5363941194A797B {1'b0}};
I13C229A5BDE90D9F920D8F4D218106DE <= 4'b0; I037773E6A298229B4A19627ABA272E81 <= 1'b0; I36FECBB048E15937DC767259CBABEDCB
<= 1'b0; end else begin I369C3845EEBC3367BADAF446789A185D <= (I84B10D95B4B5E01F827E0D4D81BF476B < 3) ? IEE94C2462F89091D3C62992327532D1E
: I88A97019335E3F57955B11E67DFFCD65 ; I13C229A5BDE90D9F920D8F4D218106DE <= (I84B10D95B4B5E01F827E0D4D81BF476B <
3) ? ((I84B10D95B4B5E01F827E0D4D81BF476B == 2) ? {IC52F3B77F7E45A74323561D6A6F6028A , {4{1'b1}}} : {{4{1'b0}}, IC52F3B77F7E45A74323561D6A6F6028A })
: {8{1'b1}}; if (IF8BC24CAD7E18C8A3A9A264889D5ECF8 ) I074FD9C5AE408613B3750B75A6125486 <= {IECBB27B02681BC7BD91D739A6D8B2975 [31:0],
I9E40C3A9F9E3CDFC05F95566701DFB02 [63:32]}; else I074FD9C5AE408613B3750B75A6125486 <= IECBB27B02681BC7BD91D739A6D8B2975 ;
end end end IF5A7A7CE92502E2DF9F0601605A38637 : begin if (I9962CDA8EE94C7BDFB23FE70815056E4 ) begin if (~IA85D446CD214F6B3CE6418205432D870 )
I26F46DF735C89C3DA76F7F404A5F650F <= 1'b1; if (I511F58CE0ACA83EE959D1BF6C4EAFA7F & ~I69B8FD7561F9CA8AAF4E50C5B2DCF850 )
begin IBFF7FD594C616C9EBAD12448149DA576 <= I71DBDE411F9CED520FD43A4EF5CBD656 ; I0C9CC98CD774EDC9DF9AB513E5A8FB57
<= 1'b1; end end else if (~IE12D7FB0707DA0B72DA8BD64B6FAEFEB ) begin if (~I45A8F29589769D54C9D702481065CB45 ) IF9A51F60DF053D68A5D57FECB5AB7ACB
<= 1'b1; if (I511F58CE0ACA83EE959D1BF6C4EAFA7F & ~IBB8FE5B389C0BD7BA64F2E05FCDC4485 ) begin I5AF6C20F3950D58007B9C0BEA7C87198
<= I71DBDE411F9CED520FD43A4EF5CBD656 ; I533559C7D3A6FC7D4A2E49A02AFC9137 <= 1'b1; end end end I5021A214EB457E909E76C621F6DD12B1
: begin IBFF7FD594C616C9EBAD12448149DA576 <= 8'b0; I0C9CC98CD774EDC9DF9AB513E5A8FB57 <= 1'b0; I26F46DF735C89C3DA76F7F404A5F650F
<= 1'b0; I5AF6C20F3950D58007B9C0BEA7C87198 <= 8'b0; I533559C7D3A6FC7D4A2E49A02AFC9137 <= 1'b0; IF9A51F60DF053D68A5D57FECB5AB7ACB
<= 1'b0; end I05E305FFF5B6CDE122F8935EE521D523 : begin I5B3BB6CF473F793585E2668A9A7136C8 <= ~I5B3BB6CF473F793585E2668A9A7136C8
| (I5B3BB6CF473F793585E2668A9A7136C8 & ~I9F4F7E2C4A4A8FB2780021EDF6E4ADEF ); end IFAC7B411ECB5421590DDAA0B7B34F238
: begin I5E1B26AB678FDA8FBEB1A0F43F21D9E4 <= I511F58CE0ACA83EE959D1BF6C4EAFA7F & ICDFF33095CB0890DA2F167B63251EC67 ;
end I248DCDE6260EE21AB43E9E1EF6D603EF : begin I5E1B26AB678FDA8FBEB1A0F43F21D9E4 <= (|I84B10D95B4B5E01F827E0D4D81BF476B )
& ~(I5E1B26AB678FDA8FBEB1A0F43F21D9E4 & ((I84B10D95B4B5E01F827E0D4D81BF476B < 3) ? 1'b1 : 1'b0)); if (IEDEC097EECBEE6B592219F6FEFFC7C2A
& (|I84B10D95B4B5E01F827E0D4D81BF476B )) begin I84B10D95B4B5E01F827E0D4D81BF476B <= (I84B10D95B4B5E01F827E0D4D81BF476B
> 1) ? I84B10D95B4B5E01F827E0D4D81BF476B - 2 : I84B10D95B4B5E01F827E0D4D81BF476B - 1; end end I6EA1237B063AFA6C82E354D0001BEF41
: begin I7FA4C54BD6B551C794EE0EA588CBD4C7 <= 1'b1; I9B8138DCE156F7C31EB5914EF01F183C <= I9119CE851F731CBC5834D0370CCA6908 [I6345C4C803C15670FB2665AEA7AA4E33 ]
| I9C46AA186B65717669AB8B1F7ED02022 ; if (I7732946249B5963DFD9C95EC611A1D2C ) if (IE655D625D2EB067AC17967E600BE5FBD )
I2C5E6805594DFF3B9EB915045ABF7575 <= {I6A62FD6104E281B8714322DB8CCB5FE3 , I18D210808E8E4FD4E19269D50B767EF6 , 10'b0,
IC4C940842A3072C3A9C40616C6A213F2 , IE8010EDEC4159FBD688A550900D0006D , I6345C4C803C15670FB2665AEA7AA4E33 , ID2A58EC9E1C805C9EA9CF0D05ACFD523 ,
1'b0, IAC85A6B0EE1F3079B60C115CB476DF06 }; else I2C5E6805594DFF3B9EB915045ABF7575 <= {I6A62FD6104E281B8714322DB8CCB5FE3 ,
I18D210808E8E4FD4E19269D50B767EF6 , 10'b0, IC4C940842A3072C3A9C40616C6A213F2 , IE8010EDEC4159FBD688A550900D0006D ,
I6345C4C803C15670FB2665AEA7AA4E33 , ID2A58EC9E1C805C9EA9CF0D05ACFD523 , 1'b0, 12'h004}; else if (IE655D625D2EB067AC17967E600BE5FBD )
I2C5E6805594DFF3B9EB915045ABF7575 <= {I85B0192F2AC4464C88E2C93352FE6696 , I18D210808E8E4FD4E19269D50B767EF6 , I30D7DB78C2B62A00872F044F1A2F39A2 [9:0],
IC4C940842A3072C3A9C40616C6A213F2 , IE8010EDEC4159FBD688A550900D0006D , I6345C4C803C15670FB2665AEA7AA4E33 , IF79BEED009A88E1D471FE1CEC77A7604 ,
1'b0, IAC85A6B0EE1F3079B60C115CB476DF06 }; else if (I511F58CE0ACA83EE959D1BF6C4EAFA7F ) I2C5E6805594DFF3B9EB915045ABF7575
<= {I6A62FD6104E281B8714322DB8CCB5FE3 , I18D210808E8E4FD4E19269D50B767EF6 , 10'b01, IC4C940842A3072C3A9C40616C6A213F2 ,
IE8010EDEC4159FBD688A550900D0006D , I6345C4C803C15670FB2665AEA7AA4E33 , IF79BEED009A88E1D471FE1CEC77A7604 , 1'b0,
12'h004}; else I2C5E6805594DFF3B9EB915045ABF7575 <= {I85B0192F2AC4464C88E2C93352FE6696 , I18D210808E8E4FD4E19269D50B767EF6 ,
10'b01, IC4C940842A3072C3A9C40616C6A213F2 , IE8010EDEC4159FBD688A550900D0006D , I6345C4C803C15670FB2665AEA7AA4E33 ,
IF79BEED009A88E1D471FE1CEC77A7604 , 1'b0, 12'h004}; I2212D954BC70C49C1F608E169DC873BC <= 1'b1; case (I11FD35FED78BCB8861FACB9A1E3A4C35 )
4'b0010, 4'b0110, 4'b1010, 4'b1110 : I54D7451A32675B2129629BC41778D6D6 <= {I83F18730E4735495B20E29C862E672F1 [6:2],
2'b01}; 4'b0100, 4'b1100 : I54D7451A32675B2129629BC41778D6D6 <= {I83F18730E4735495B20E29C862E672F1 [6:2], 2'b10};
4'b1000 : I54D7451A32675B2129629BC41778D6D6 <= {I83F18730E4735495B20E29C862E672F1 [6:2], 2'b11}; default I54D7451A32675B2129629BC41778D6D6
<= I83F18730E4735495B20E29C862E672F1 [6:0]; endcase end I070181DB2ED3EDD3633DB4E93B8E42A5 : begin if (IE655D625D2EB067AC17967E600BE5FBD )
I2C5E6805594DFF3B9EB915045ABF7575 <= {IB9A23596C80981B9B1CF7E12A76E71AC , I288715DFB3893A064D51571152559F12 , I86B9557FA0123B8105E34300F4FCD447 ,
I539C1D01FC349447001EB93E17D37611 , 1'b0, I54D7451A32675B2129629BC41778D6D6 , {32{1'b0}}}; else I2C5E6805594DFF3B9EB915045ABF7575
<= {IB9A23596C80981B9B1CF7E12A76E71AC , I288715DFB3893A064D51571152559F12 , I86B9557FA0123B8105E34300F4FCD447 ,
I539C1D01FC349447001EB93E17D37611 , 1'b0, 7'b0, {32{1'b0}}}; I893DF0D582AF0617B44879E65C202360 <= I7732946249B5963DFD9C95EC611A1D2C
| I511F58CE0ACA83EE959D1BF6C4EAFA7F ; I2212D954BC70C49C1F608E169DC873BC <= I7732946249B5963DFD9C95EC611A1D2C | I511F58CE0ACA83EE959D1BF6C4EAFA7F ;
end I2263EE3B1CDD9957F685B729A9639643 : begin IF8BC24CAD7E18C8A3A9A264889D5ECF8 <= ~I54D7451A32675B2129629BC41778D6D6 [2];
I893DF0D582AF0617B44879E65C202360 <= 1'b0; I2212D954BC70C49C1F608E169DC873BC <= 1'b0; if (I511F58CE0ACA83EE959D1BF6C4EAFA7F )
I2C5E6805594DFF3B9EB915045ABF7575 <= {64{1'b0}}; end endcase end end endmodule 
 module I4A464F8B941F768B40777E11E08CF0DE # (parameter I7292F55C07BFD7FB8A60D29FFC186275 = 32, parameter IDB9D60794264C5F8E5363941194A797B
= 3, parameter ID7C7F9F2E39BEBEE2ACFA8040034E48D = 24 ) ( input wire ICCFB0F435B37370076102F325BC08D20 , input wire
I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire IAB4F3026BD4F2760154E70C5BC0FE751 , input wire [I7292F55C07BFD7FB8A60D29FFC186275
- 1:0] ID8E639B3434FEAB4D1CA5AF230310D49 , input wire IC43B0BCCD0A723BBF62FF7B9D230C3F8 , input wire I122CA37F449B813A5F0CAF8BC20EE9EA ,
input wire IFD5EF944B5EFFB20EE3422B3D79A2BF4 , input wire IB7C0B3EE4A87531F21610094A69146A7 , input wire IF87783FDF111A8E49EAC36F1DDFCBA80 ,
input wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] IF9D5978BE23690B1D4D13EF2AD676C6F , input wire [ID7C7F9F2E39BEBEE2ACFA8040034E48D
- 1:0] IDC6EA54AB52AEAD439CEF7521615AE1B , input wire [2:0] I6ED49B5BED4BA586759FFDCC7B3B7FF8 , input wire [IDB9D60794264C5F8E5363941194A797B
- 1:0] I8E2F7CF6E50B95A483351A1836EB23AC , input wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] I506D2FCB600E0189274870B654E65B64 ,
input wire I141300E29D7EF4A0D8B71CB7469A7B90 , input wire I9AF8DD3F367CE82DF45437DB546EAAD3 , input wire [10:0]
I42D281FF99DC79A9AD9E7DF0AEB073A7 , input wire [3:0] I3068B33EE97A971AE7F0CF17705AA6DC , input wire [3:0] IFCBA19703D55B4610B3F4174C5B8833A ,
input wire IC3CC91D317012C130AC9E2A126F71C64 , output wire ID8C32104758E11D83079BB9AEE0C35DB , output wire IC91681A00788ED1B6C6956634033ED38 ,
output wire I7114A89BF31DB18ED21FF0608A9BF50A , output wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] IB2B35E1DF060E7BC2B7E414954F6FA34 ,
output wire [ID7C7F9F2E39BEBEE2ACFA8040034E48D - 1:0] I561BE0F01153FC1AADDEB08B34B545B6 , output wire [1:0] IB86AF6EBEEA3CE1BF22AE1AF7CC8481F ,
output wire [2:0] I94E3D00BBC13BF182097A25D63288C2C , output wire [IDB9D60794264C5F8E5363941194A797B - 1:0] I8B25F4450817FC10E1E3DC6B500C9F5A ,
output wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] I26C902CE18647F75561AD003E260B048 , output wire [3:0] IA5CEBFC654EDCA4107594F388D5BC88A ,
output wire I27627079DD78A85D26D85DC0C53D835F , output wire I0205131FB84BB0F9F8AD5CC00E5E861D , output wire IDA581E8478C8224118EF4E6B8EE8DDFE ,
output wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] IA36C0DD0DE88B03FA61EF35103D22DF0 ); `include "wishbone_utils.v"
 localparam IFD36C31411244EF5908C439ABA23D673 = 3'b000, IE42F0B27BC424D7A06FC837E3293B736 = 3'b001, I1CFF64FE635B8A5E53C413D36FBCCCB2
= 3'b010, I9D1C0AC088DEB1CAC7C2753E2CBDE708 = 3'b011, I8EB8B007E61CF9BBAD642C3B9D452755 = 3'b100, IAA47CC78E75AE27D93BDEFEEAA1D9FE0
= 3'b101, I8C5E7A65ED8A08585AFDA3F064E91620 = 3'b110;  reg I83C48096FC314C76A39446D6CEC94A5E ; reg I3B7C6E5488B3FB1985C6E71FB483FEAC ;
reg [11:0] IFC80E6824CDF033E77AC2726508CCAF2 ; reg [ID7C7F9F2E39BEBEE2ACFA8040034E48D - 1:0] IC7779D4175ADF3F75C21392F9E824B6D ;
reg [1:0] IA6B00370F90E5BFE7B5D8852390CF107 ; reg [2:0] I369C3845EEBC3367BADAF446789A185D ; reg [IDB9D60794264C5F8E5363941194A797B
- 1:0] ID564A30F71C7C1B827BA57264E89B21D ; reg [2:0] I15BDB8EF2F82D399EEAB37F26106A134 ; reg [2:0] I611306DB4017E4CC74DC60EB7716CFC8 ;
reg [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] I3EAE45CFB73C88FE02CA1913C5C393B0 ; reg [3:0] I13C229A5BDE90D9F920D8F4D218106DE ;
reg I037773E6A298229B4A19627ABA272E81 ; reg [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] IE52F11681C095BD0BF82CB1F94B17953 ;
reg I36FECBB048E15937DC767259CBABEDCB ; reg [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] I185849505AD09166EC514C856BD76D16 ;
reg I744748C802A4982FBAC6677930DA7B4E ; reg I2D1C4F8EF2C236DEEDB8729F3B943A14 ; reg I077A22296F5A2EAC26F7E1C101A6DD66 ;
reg IFE5A0EABD9C5876584C2797DD70F1C53 ; reg [ID7C7F9F2E39BEBEE2ACFA8040034E48D - 1:0] IBB9F765CF2FE61A77D4144021BAD1FF3 ;
reg [11:0] I8244A0A6CFBB12A29C0A59DBB4FC13EE ; reg [IDB9D60794264C5F8E5363941194A797B - 1:0] I2A11E8CA4C8D03C39CA9F863A29AC507 ;
reg IFD5BC87AA0B9E0C4586F686D5FDF1E99 ; reg I3BFFD10A33B9292FB529E91CBF53786E ; reg [3:0] I31DFC7DC35DC851D2F9F524A08DCA457 ;
reg [3:0] I9D1E56BC71C6D6CEB6D98E56F8B5C157 ; reg I92697AA5627C77767A135FE38B5E0E73 ; wire IF2AFEE13983D94D5364425E9CE96BD48 ;
wire ID408E2DFA2D752FEF4954B0FB0BED658 ; wire I9B39837C897B4C3F93D215848CAA866E ; wire I3198775D45BDCB2F4B3A4E26EEB19AF8 ;
wire I6F92245E15C786DD863084D65306C438 ;  assign ID8C32104758E11D83079BB9AEE0C35DB = I83C48096FC314C76A39446D6CEC94A5E ;
assign IC91681A00788ED1B6C6956634033ED38 = I3B7C6E5488B3FB1985C6E71FB483FEAC | IF2AFEE13983D94D5364425E9CE96BD48 ;
assign I7114A89BF31DB18ED21FF0608A9BF50A = ID408E2DFA2D752FEF4954B0FB0BED658 ; assign IB2B35E1DF060E7BC2B7E414954F6FA34
= (I077A22296F5A2EAC26F7E1C101A6DD66 & ~I92697AA5627C77767A135FE38B5E0E73 ) ? I3EAE45CFB73C88FE02CA1913C5C393B0
: I506D2FCB600E0189274870B654E65B64 ; assign I561BE0F01153FC1AADDEB08B34B545B6 = IC7779D4175ADF3F75C21392F9E824B6D ;
assign IB86AF6EBEEA3CE1BF22AE1AF7CC8481F = IA6B00370F90E5BFE7B5D8852390CF107 ; assign I94E3D00BBC13BF182097A25D63288C2C
= I369C3845EEBC3367BADAF446789A185D ; assign I8B25F4450817FC10E1E3DC6B500C9F5A = ID564A30F71C7C1B827BA57264E89B21D ;
assign I26C902CE18647F75561AD003E260B048 = IE52F11681C095BD0BF82CB1F94B17953 ; assign IA5CEBFC654EDCA4107594F388D5BC88A
= I13C229A5BDE90D9F920D8F4D218106DE ; assign I27627079DD78A85D26D85DC0C53D835F = I037773E6A298229B4A19627ABA272E81 ;
assign I0205131FB84BB0F9F8AD5CC00E5E861D = I36FECBB048E15937DC767259CBABEDCB ; assign IDA581E8478C8224118EF4E6B8EE8DDFE
= I9B39837C897B4C3F93D215848CAA866E ; assign IA36C0DD0DE88B03FA61EF35103D22DF0 = (IFE5A0EABD9C5876584C2797DD70F1C53 )
? I185849505AD09166EC514C856BD76D16 : {I7292F55C07BFD7FB8A60D29FFC186275 {1'b0}};  assign IF2AFEE13983D94D5364425E9CE96BD48
= I077A22296F5A2EAC26F7E1C101A6DD66 & I92697AA5627C77767A135FE38B5E0E73 & I141300E29D7EF4A0D8B71CB7469A7B90 & I9B39837C897B4C3F93D215848CAA866E ;
assign ID408E2DFA2D752FEF4954B0FB0BED658 = ((I077A22296F5A2EAC26F7E1C101A6DD66 == 1'b1) && (I92697AA5627C77767A135FE38B5E0E73
== 1'b1)) ? ((|ID564A30F71C7C1B827BA57264E89B21D ) & ~IF87783FDF111A8E49EAC36F1DDFCBA80 ) : 1'b0; assign I9B39837C897B4C3F93D215848CAA866E
= (I077A22296F5A2EAC26F7E1C101A6DD66 ) ? ((I92697AA5627C77767A135FE38B5E0E73 ) ? (~(I122CA37F449B813A5F0CAF8BC20EE9EA
| I2D1C4F8EF2C236DEEDB8729F3B943A14 )) : I744748C802A4982FBAC6677930DA7B4E ) : 1'b0; assign I3198775D45BDCB2F4B3A4E26EEB19AF8
= (I6ED49B5BED4BA586759FFDCC7B3B7FF8 == IEE94C2462F89091D3C62992327532D1E ) ? (I141300E29D7EF4A0D8B71CB7469A7B90
& I9B39837C897B4C3F93D215848CAA866E ) : 1'b0; assign I6F92245E15C786DD863084D65306C438 = (I141300E29D7EF4A0D8B71CB7469A7B90
& (|I8E2F7CF6E50B95A483351A1836EB23AC ) & ~IC3CC91D317012C130AC9E2A126F71C64 ) | ((|I8E2F7CF6E50B95A483351A1836EB23AC )
& IC3CC91D317012C130AC9E2A126F71C64 );  always @(*) begin I611306DB4017E4CC74DC60EB7716CFC8 = I15BDB8EF2F82D399EEAB37F26106A134 ;
case (I15BDB8EF2F82D399EEAB37F26106A134 ) IFD36C31411244EF5908C439ABA23D673 : begin if (I6F92245E15C786DD863084D65306C438 )
I611306DB4017E4CC74DC60EB7716CFC8 = IE42F0B27BC424D7A06FC837E3293B736 ; end IE42F0B27BC424D7A06FC837E3293B736 :
begin if (I92697AA5627C77767A135FE38B5E0E73 ) begin if (IC43B0BCCD0A723BBF62FF7B9D230C3F8 == 1'b0) I611306DB4017E4CC74DC60EB7716CFC8
= I1CFF64FE635B8A5E53C413D36FBCCCB2 ; end else begin if (IC43B0BCCD0A723BBF62FF7B9D230C3F8 == 1'b1) I611306DB4017E4CC74DC60EB7716CFC8
= I1CFF64FE635B8A5E53C413D36FBCCCB2 ; end end I1CFF64FE635B8A5E53C413D36FBCCCB2 : begin if (I92697AA5627C77767A135FE38B5E0E73 )
I611306DB4017E4CC74DC60EB7716CFC8 = I9D1C0AC088DEB1CAC7C2753E2CBDE708 ; else I611306DB4017E4CC74DC60EB7716CFC8 =
I8EB8B007E61CF9BBAD642C3B9D452755 ; end I9D1C0AC088DEB1CAC7C2753E2CBDE708 : begin if (IB7C0B3EE4A87531F21610094A69146A7
== 1'b1) I611306DB4017E4CC74DC60EB7716CFC8 = IAA47CC78E75AE27D93BDEFEEAA1D9FE0 ; end I8EB8B007E61CF9BBAD642C3B9D452755
: begin if (I3BFFD10A33B9292FB529E91CBF53786E & I037773E6A298229B4A19627ABA272E81 & IF87783FDF111A8E49EAC36F1DDFCBA80 )
I611306DB4017E4CC74DC60EB7716CFC8 = I8C5E7A65ED8A08585AFDA3F064E91620 ; end IAA47CC78E75AE27D93BDEFEEAA1D9FE0 :
begin if (I3BFFD10A33B9292FB529E91CBF53786E & I037773E6A298229B4A19627ABA272E81 & IF87783FDF111A8E49EAC36F1DDFCBA80 )
I611306DB4017E4CC74DC60EB7716CFC8 = IFD36C31411244EF5908C439ABA23D673 ; end I8C5E7A65ED8A08585AFDA3F064E91620 :
begin if (I3198775D45BDCB2F4B3A4E26EEB19AF8 ) I611306DB4017E4CC74DC60EB7716CFC8 = IFD36C31411244EF5908C439ABA23D673 ;
end endcase end  always @(posedge ICCFB0F435B37370076102F325BC08D20 or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 )
if (~I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin I83C48096FC314C76A39446D6CEC94A5E <= 1'b0; I3B7C6E5488B3FB1985C6E71FB483FEAC
<= 1'b0; IFC80E6824CDF033E77AC2726508CCAF2 <= 11'b0; IC7779D4175ADF3F75C21392F9E824B6D <= {ID7C7F9F2E39BEBEE2ACFA8040034E48D {1'b0}};
IA6B00370F90E5BFE7B5D8852390CF107 <= {2{1'b0}}; I369C3845EEBC3367BADAF446789A185D <= {3{1'b0}}; ID564A30F71C7C1B827BA57264E89B21D
<= {IDB9D60794264C5F8E5363941194A797B {1'b0}}; I15BDB8EF2F82D399EEAB37F26106A134 <= IFD36C31411244EF5908C439ABA23D673 ;
I3EAE45CFB73C88FE02CA1913C5C393B0 <= {I7292F55C07BFD7FB8A60D29FFC186275 {1'b0}}; I13C229A5BDE90D9F920D8F4D218106DE
<= {4{1'b0}}; I037773E6A298229B4A19627ABA272E81 <= 1'b0; IE52F11681C095BD0BF82CB1F94B17953 <= {I7292F55C07BFD7FB8A60D29FFC186275 {1'b0}};
I36FECBB048E15937DC767259CBABEDCB <= 1'b0; I185849505AD09166EC514C856BD76D16 <= {I7292F55C07BFD7FB8A60D29FFC186275 {1'b0}};
I744748C802A4982FBAC6677930DA7B4E <= 1'b0; I2D1C4F8EF2C236DEEDB8729F3B943A14 <= 1'b0; I077A22296F5A2EAC26F7E1C101A6DD66
<= 1'b0; IFE5A0EABD9C5876584C2797DD70F1C53 <= 1'b0; IBB9F765CF2FE61A77D4144021BAD1FF3 <= {ID7C7F9F2E39BEBEE2ACFA8040034E48D {1'b0}};
I8244A0A6CFBB12A29C0A59DBB4FC13EE <= {11{1'b0}}; I2A11E8CA4C8D03C39CA9F863A29AC507 <= {IDB9D60794264C5F8E5363941194A797B {1'b0}};
IFD5BC87AA0B9E0C4586F686D5FDF1E99 <= 1'b0; I3BFFD10A33B9292FB529E91CBF53786E <= 1'b0; I31DFC7DC35DC851D2F9F524A08DCA457
<= {4{1'b0}}; I9D1E56BC71C6D6CEB6D98E56F8B5C157 <= {4{1'b0}}; I92697AA5627C77767A135FE38B5E0E73 <= 1'b0; end else
begin I83C48096FC314C76A39446D6CEC94A5E <= (IFC80E6824CDF033E77AC2726508CCAF2 > 0) ? ((~I92697AA5627C77767A135FE38B5E0E73
& ~IC43B0BCCD0A723BBF62FF7B9D230C3F8 & ~(I83C48096FC314C76A39446D6CEC94A5E & IFD5EF944B5EFFB20EE3422B3D79A2BF4 ))
| (I92697AA5627C77767A135FE38B5E0E73 & ~IC43B0BCCD0A723BBF62FF7B9D230C3F8 & ~(I83C48096FC314C76A39446D6CEC94A5E
& IFD5EF944B5EFFB20EE3422B3D79A2BF4 ) & ~((|ID564A30F71C7C1B827BA57264E89B21D ) & ~IF87783FDF111A8E49EAC36F1DDFCBA80 )))
: 1'b0; I3B7C6E5488B3FB1985C6E71FB483FEAC <= 1'b0; I15BDB8EF2F82D399EEAB37F26106A134 <= I611306DB4017E4CC74DC60EB7716CFC8 ;
I185849505AD09166EC514C856BD76D16 <= (I92697AA5627C77767A135FE38B5E0E73 == 1'b0) ? ID8E639B3434FEAB4D1CA5AF230310D49
: {I7292F55C07BFD7FB8A60D29FFC186275 {1'b0}}; I744748C802A4982FBAC6677930DA7B4E <= IB7C0B3EE4A87531F21610094A69146A7
& ~I92697AA5627C77767A135FE38B5E0E73 ; I2D1C4F8EF2C236DEEDB8729F3B943A14 <= (I15BDB8EF2F82D399EEAB37F26106A134 ==
IFD36C31411244EF5908C439ABA23D673 ) ? 1'b0 : (I2D1C4F8EF2C236DEEDB8729F3B943A14 | (I077A22296F5A2EAC26F7E1C101A6DD66
& I3198775D45BDCB2F4B3A4E26EEB19AF8 )); if (IFC80E6824CDF033E77AC2726508CCAF2 > 0) begin if (I83C48096FC314C76A39446D6CEC94A5E
& ~ID408E2DFA2D752FEF4954B0FB0BED658 ) IFC80E6824CDF033E77AC2726508CCAF2 <= IFC80E6824CDF033E77AC2726508CCAF2 -
1; end case (I15BDB8EF2F82D399EEAB37F26106A134 ) IFD36C31411244EF5908C439ABA23D673 : begin if (I6F92245E15C786DD863084D65306C438 )
begin I077A22296F5A2EAC26F7E1C101A6DD66 <= 1'b1; IFE5A0EABD9C5876584C2797DD70F1C53 <= ~IC3CC91D317012C130AC9E2A126F71C64 ;
IBB9F765CF2FE61A77D4144021BAD1FF3 <= IDC6EA54AB52AEAD439CEF7521615AE1B ; I8244A0A6CFBB12A29C0A59DBB4FC13EE <= I42D281FF99DC79A9AD9E7DF0AEB073A7 ;
I2A11E8CA4C8D03C39CA9F863A29AC507 <= I8E2F7CF6E50B95A483351A1836EB23AC ; I31DFC7DC35DC851D2F9F524A08DCA457 <= I3068B33EE97A971AE7F0CF17705AA6DC ;
I9D1E56BC71C6D6CEB6D98E56F8B5C157 <= IFCBA19703D55B4610B3F4174C5B8833A ; I92697AA5627C77767A135FE38B5E0E73 <= IC3CC91D317012C130AC9E2A126F71C64 ;
end end IE42F0B27BC424D7A06FC837E3293B736 : begin IFD5BC87AA0B9E0C4586F686D5FDF1E99 <= (I8244A0A6CFBB12A29C0A59DBB4FC13EE
== 2) ? 1'b1 : 1'b0; I3BFFD10A33B9292FB529E91CBF53786E <= (I8244A0A6CFBB12A29C0A59DBB4FC13EE == 1) ? 1'b1 : 1'b0;
end I1CFF64FE635B8A5E53C413D36FBCCCB2 : begin IFC80E6824CDF033E77AC2726508CCAF2 <= I8244A0A6CFBB12A29C0A59DBB4FC13EE ;
if (~I92697AA5627C77767A135FE38B5E0E73 ) begin IC7779D4175ADF3F75C21392F9E824B6D <= IBB9F765CF2FE61A77D4144021BAD1FF3 ;
IA6B00370F90E5BFE7B5D8852390CF107 <= 2'b0; I369C3845EEBC3367BADAF446789A185D <= (I3BFFD10A33B9292FB529E91CBF53786E )
? IEE94C2462F89091D3C62992327532D1E : I88A97019335E3F57955B11E67DFFCD65 ; ID564A30F71C7C1B827BA57264E89B21D <= I2A11E8CA4C8D03C39CA9F863A29AC507 ;
I13C229A5BDE90D9F920D8F4D218106DE <= I31DFC7DC35DC851D2F9F524A08DCA457 ; I037773E6A298229B4A19627ABA272E81 <= 1'b1;
IE52F11681C095BD0BF82CB1F94B17953 <= {I7292F55C07BFD7FB8A60D29FFC186275 {1'b0}}; I36FECBB048E15937DC767259CBABEDCB
<= 1'b0; end end I9D1C0AC088DEB1CAC7C2753E2CBDE708 : begin if (IB7C0B3EE4A87531F21610094A69146A7 == 1'b1) begin
IC7779D4175ADF3F75C21392F9E824B6D <= IBB9F765CF2FE61A77D4144021BAD1FF3 ; IA6B00370F90E5BFE7B5D8852390CF107 <= 2'b0;
I369C3845EEBC3367BADAF446789A185D <= (I3BFFD10A33B9292FB529E91CBF53786E ) ? IEE94C2462F89091D3C62992327532D1E :
I88A97019335E3F57955B11E67DFFCD65 ; ID564A30F71C7C1B827BA57264E89B21D <= I2A11E8CA4C8D03C39CA9F863A29AC507 ; I13C229A5BDE90D9F920D8F4D218106DE
<= I31DFC7DC35DC851D2F9F524A08DCA457 ; I037773E6A298229B4A19627ABA272E81 <= 1'b1; IE52F11681C095BD0BF82CB1F94B17953
<= ID8E639B3434FEAB4D1CA5AF230310D49 ; I36FECBB048E15937DC767259CBABEDCB <= 1'b1; end end I8EB8B007E61CF9BBAD642C3B9D452755
: begin if (I037773E6A298229B4A19627ABA272E81 & IF87783FDF111A8E49EAC36F1DDFCBA80 ) begin I3B7C6E5488B3FB1985C6E71FB483FEAC
<= 1'b1; I8244A0A6CFBB12A29C0A59DBB4FC13EE <= I8244A0A6CFBB12A29C0A59DBB4FC13EE - 1; IFD5BC87AA0B9E0C4586F686D5FDF1E99
<= (I8244A0A6CFBB12A29C0A59DBB4FC13EE == 3) ? 1'b1 : 1'b0; I3BFFD10A33B9292FB529E91CBF53786E <= (I8244A0A6CFBB12A29C0A59DBB4FC13EE
== 2) ? 1'b1 : 1'b0; I3EAE45CFB73C88FE02CA1913C5C393B0 <= IF9D5978BE23690B1D4D13EF2AD676C6F ; if (I3BFFD10A33B9292FB529E91CBF53786E )
begin IC7779D4175ADF3F75C21392F9E824B6D <= {ID7C7F9F2E39BEBEE2ACFA8040034E48D {1'b0}}; IA6B00370F90E5BFE7B5D8852390CF107
<= {2{1'b0}}; I369C3845EEBC3367BADAF446789A185D <= {3{1'b0}}; ID564A30F71C7C1B827BA57264E89B21D <= {IDB9D60794264C5F8E5363941194A797B {1'b0}};
I13C229A5BDE90D9F920D8F4D218106DE <= {4{1'b0}}; I037773E6A298229B4A19627ABA272E81 <= 1'b0; IE52F11681C095BD0BF82CB1F94B17953
<= {I7292F55C07BFD7FB8A60D29FFC186275 {1'b0}}; I36FECBB048E15937DC767259CBABEDCB <= 1'b0; end else begin IC7779D4175ADF3F75C21392F9E824B6D
<= IC7779D4175ADF3F75C21392F9E824B6D + 4; I369C3845EEBC3367BADAF446789A185D <= (IFD5BC87AA0B9E0C4586F686D5FDF1E99 )
? IEE94C2462F89091D3C62992327532D1E : I88A97019335E3F57955B11E67DFFCD65 ; I13C229A5BDE90D9F920D8F4D218106DE <= (IFD5BC87AA0B9E0C4586F686D5FDF1E99 )
? I9D1E56BC71C6D6CEB6D98E56F8B5C157 : {4{1'b1}}; I037773E6A298229B4A19627ABA272E81 <= ~IAB4F3026BD4F2760154E70C5BC0FE751 ;
end end else begin I037773E6A298229B4A19627ABA272E81 <= I037773E6A298229B4A19627ABA272E81 | (~I037773E6A298229B4A19627ABA272E81
& ~IAB4F3026BD4F2760154E70C5BC0FE751 ); end end IAA47CC78E75AE27D93BDEFEEAA1D9FE0 : begin if (I037773E6A298229B4A19627ABA272E81
& IF87783FDF111A8E49EAC36F1DDFCBA80 ) begin I8244A0A6CFBB12A29C0A59DBB4FC13EE <= I8244A0A6CFBB12A29C0A59DBB4FC13EE
- 1; IFD5BC87AA0B9E0C4586F686D5FDF1E99 <= (I8244A0A6CFBB12A29C0A59DBB4FC13EE == 3) ? 1'b1 : 1'b0; I3BFFD10A33B9292FB529E91CBF53786E
<= (I8244A0A6CFBB12A29C0A59DBB4FC13EE == 2) ? 1'b1 : 1'b0; if (I3BFFD10A33B9292FB529E91CBF53786E ) begin IC7779D4175ADF3F75C21392F9E824B6D
<= {ID7C7F9F2E39BEBEE2ACFA8040034E48D {1'b0}}; IA6B00370F90E5BFE7B5D8852390CF107 <= {2{1'b0}}; I369C3845EEBC3367BADAF446789A185D
<= {3{1'b0}}; ID564A30F71C7C1B827BA57264E89B21D <= {IDB9D60794264C5F8E5363941194A797B {1'b0}}; I13C229A5BDE90D9F920D8F4D218106DE
<= {4{1'b0}}; I037773E6A298229B4A19627ABA272E81 <= 1'b0; IE52F11681C095BD0BF82CB1F94B17953 <= {I7292F55C07BFD7FB8A60D29FFC186275 {1'b0}};
I36FECBB048E15937DC767259CBABEDCB <= 1'b0; I077A22296F5A2EAC26F7E1C101A6DD66 <= 1'b0; IFE5A0EABD9C5876584C2797DD70F1C53
<= 1'b0; end else begin IC7779D4175ADF3F75C21392F9E824B6D <= IC7779D4175ADF3F75C21392F9E824B6D + 4; I369C3845EEBC3367BADAF446789A185D
<= (IFD5BC87AA0B9E0C4586F686D5FDF1E99 ) ? IEE94C2462F89091D3C62992327532D1E : I88A97019335E3F57955B11E67DFFCD65 ;
I13C229A5BDE90D9F920D8F4D218106DE <= (IFD5BC87AA0B9E0C4586F686D5FDF1E99 ) ? I9D1E56BC71C6D6CEB6D98E56F8B5C157 :
{4{1'b1}}; I037773E6A298229B4A19627ABA272E81 <= IB7C0B3EE4A87531F21610094A69146A7 ; IE52F11681C095BD0BF82CB1F94B17953
<= (IB7C0B3EE4A87531F21610094A69146A7 == 1'b1) ? ID8E639B3434FEAB4D1CA5AF230310D49 : IE52F11681C095BD0BF82CB1F94B17953 ;
end end else begin I037773E6A298229B4A19627ABA272E81 <= I037773E6A298229B4A19627ABA272E81 | IB7C0B3EE4A87531F21610094A69146A7 ;
IE52F11681C095BD0BF82CB1F94B17953 <= (IB7C0B3EE4A87531F21610094A69146A7 & ~I037773E6A298229B4A19627ABA272E81 ) ?
ID8E639B3434FEAB4D1CA5AF230310D49 : IE52F11681C095BD0BF82CB1F94B17953 ; end end I8C5E7A65ED8A08585AFDA3F064E91620
: begin I077A22296F5A2EAC26F7E1C101A6DD66 <= ~I3198775D45BDCB2F4B3A4E26EEB19AF8 ; IFE5A0EABD9C5876584C2797DD70F1C53
<= IFE5A0EABD9C5876584C2797DD70F1C53 & ~I3198775D45BDCB2F4B3A4E26EEB19AF8 ; end endcase end endmodule 
  module I35D01845B6D15D59E4E7B95EDE6F3368 #( parameter I7292F55C07BFD7FB8A60D29FFC186275 = 32, parameter IB71844FFA3AB85FEF45EAB4D35395752
= 512, parameter IDB9D60794264C5F8E5363941194A797B = 3, parameter I66C185998F46A7148163982E39BCD296 = "ecp3", parameter
ID7C7F9F2E39BEBEE2ACFA8040034E48D = 24 ) ( input wire ICCFB0F435B37370076102F325BC08D20 , input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 ,
input wire IF87783FDF111A8E49EAC36F1DDFCBA80 , input wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] IF9D5978BE23690B1D4D13EF2AD676C6F ,
input wire [ID7C7F9F2E39BEBEE2ACFA8040034E48D - 1:0] IDC6EA54AB52AEAD439CEF7521615AE1B , input wire [2:0] I6ED49B5BED4BA586759FFDCC7B3B7FF8 ,
input wire [IDB9D60794264C5F8E5363941194A797B - 1:0] I8E2F7CF6E50B95A483351A1836EB23AC , input wire [I7292F55C07BFD7FB8A60D29FFC186275
- 1:0] I506D2FCB600E0189274870B654E65B64 , input wire I141300E29D7EF4A0D8B71CB7469A7B90 , input wire I9AF8DD3F367CE82DF45437DB546EAAD3 ,
input wire [10:0] I42D281FF99DC79A9AD9E7DF0AEB073A7 , input wire [3:0] I3068B33EE97A971AE7F0CF17705AA6DC , input
wire [3:0] IFCBA19703D55B4610B3F4174C5B8833A , input wire IC3CC91D317012C130AC9E2A126F71C64 , output wire [ID7C7F9F2E39BEBEE2ACFA8040034E48D
- 1:0] I561BE0F01153FC1AADDEB08B34B545B6 , output wire [1:0] IB86AF6EBEEA3CE1BF22AE1AF7CC8481F , output wire [2:0]
I94E3D00BBC13BF182097A25D63288C2C , output wire [IDB9D60794264C5F8E5363941194A797B - 1:0] I8B25F4450817FC10E1E3DC6B500C9F5A ,
output wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] I26C902CE18647F75561AD003E260B048 , output wire [3:0] IA5CEBFC654EDCA4107594F388D5BC88A ,
output wire I27627079DD78A85D26D85DC0C53D835F , output wire I0205131FB84BB0F9F8AD5CC00E5E861D , output wire IDA581E8478C8224118EF4E6B8EE8DDFE ,
output wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] IA36C0DD0DE88B03FA61EF35103D22DF0 );  localparam integer I36A1B4EB5B5564A6ED7EA4D42856EFB4
= $clog2(IB71844FFA3AB85FEF45EAB4D35395752 ); localparam integer I2F8DC10449A1F24468235753BBC3B988 = $clog2(IB71844FFA3AB85FEF45EAB4D35395752
+ 1); localparam integer IF35F7B506981B2912E2486B227CB8871 = I7292F55C07BFD7FB8A60D29FFC186275 ;  wire I4AE98FF3DA4D5A5EE68F8A14D9D781F4 ;
wire [I36A1B4EB5B5564A6ED7EA4D42856EFB4 - 1:0] IC2A6ECC367E2C82B97E73A57A8A79E1A ; wire I60B15FF62AA99717C8B7DA7D6912D281 ;
wire ICB86B570A185B89048AE76A09444BA41 ; wire IA6BBDC90BCC6EF2E35BFA8D709343BF3 ; wire [I36A1B4EB5B5564A6ED7EA4D42856EFB4
- 1:0] I5631F39935597168A2C9D3656C66CB5C ; wire I0E620501249C5CFBF447631D04D33715 ; wire I25891FD4BF8EA7F9051CE324A21ED31E ;
wire I366EB0B781FD462E1BDC374519E76C20 ; wire [IF35F7B506981B2912E2486B227CB8871 - 1:0] I2CA1A324143051A0AFDEFB54659C657C ;
wire I76EFAFF6D4391A79F5CD2CA7904431E8 ; wire IAFB0D72A35BE81312B83F6EC64D8ECF4 ; wire I9AC67CC0D048C17AC2F808C22F4DEE6F ;
wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] IFD939E5BC1AA3DCE57CCDC18CA4F72A8 ; wire [ID7C7F9F2E39BEBEE2ACFA8040034E48D
- 1:0] I6EFB980269078EDFE25D9139188C0357 ; wire [1:0] ID6BA376F6FDCA561D55334C951D81896 ; wire [2:0] I1261C037D95D7AC9FB55409369EA711E ;
wire [IDB9D60794264C5F8E5363941194A797B - 1:0] IAB4361F44053B3532F19F9BCB33E265F ; wire [I7292F55C07BFD7FB8A60D29FFC186275
- 1:0] I51F8ACA4F6E2B0688214E337318D090C ; wire [3:0] IAC7F9C0E3110EC41B40E14F4AFDB4D41 ; wire I3645064ACD6F902F18DE49FBB6F7350B ;
wire I64F37E01600233FCC804B26C0900CDE5 ; wire ICA81D2D21EB4C7C4D7C6096277C9D15A ; wire [I7292F55C07BFD7FB8A60D29FFC186275
- 1:0] I200E0F93328C05371EF92973FC08E636 ; wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] I081545483B2E87A5F84E4E80F8AD87A7 ;
wire IE664D85E83E89DA36250C2ADD2CC9541 ; wire IE43DA634E45C0D88369455568042AF37 ;  assign I561BE0F01153FC1AADDEB08B34B545B6
= I6EFB980269078EDFE25D9139188C0357 ; assign IB86AF6EBEEA3CE1BF22AE1AF7CC8481F = ID6BA376F6FDCA561D55334C951D81896 ;
assign I94E3D00BBC13BF182097A25D63288C2C = I1261C037D95D7AC9FB55409369EA711E ; assign I8B25F4450817FC10E1E3DC6B500C9F5A
= IAB4361F44053B3532F19F9BCB33E265F ; assign I26C902CE18647F75561AD003E260B048 = I51F8ACA4F6E2B0688214E337318D090C ;
assign IA5CEBFC654EDCA4107594F388D5BC88A = IAC7F9C0E3110EC41B40E14F4AFDB4D41 ; assign I27627079DD78A85D26D85DC0C53D835F
= I3645064ACD6F902F18DE49FBB6F7350B ; assign I0205131FB84BB0F9F8AD5CC00E5E861D = I64F37E01600233FCC804B26C0900CDE5 ;
assign IDA581E8478C8224118EF4E6B8EE8DDFE = ICA81D2D21EB4C7C4D7C6096277C9D15A ; assign IA36C0DD0DE88B03FA61EF35103D22DF0
= I200E0F93328C05371EF92973FC08E636 ;  assign I4AE98FF3DA4D5A5EE68F8A14D9D781F4 = ~I9ED2A9117D3AEAF54CBA7AD69083BCB7 ;
 IF50ADBFC5F4E76B680AD98E97599279A #( .I5D7F61632782AFE440ADE65900D53412 (2), .I61D0345D311EC6FFC08DDDECE5F6127A
(IB71844FFA3AB85FEF45EAB4D35395752 ) ) IB420C4D1279F971E867FA537CA4D6E82 ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ),
.I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .IC79EC9A9F373F4B71374BDF6EDD31DE6 (1'b0),
.ID8853B025150C80EE45BBA98E5BEA3A8 (IE664D85E83E89DA36250C2ADD2CC9541 ), .I22B24791BA0E7AA2C686B1B2D776C636 (IAFB0D72A35BE81312B83F6EC64D8ECF4 ),
.I79D313D86841E5141E7629EA606D7AE9 (IC2A6ECC367E2C82B97E73A57A8A79E1A ), .I11CEFC90537A67CD1FF01400245362F2 ( ),
.ID7FCE45A65ADDB17F91F73A1B506BB5B ( ), .I8BB939FF2AFDE7B2A1E480DCB61CE354 (I60B15FF62AA99717C8B7DA7D6912D281 ),
.I41C63F948E534C7ED9F2471A44C922B2 (ICB86B570A185B89048AE76A09444BA41 ), .I585F74DE05DD9C1C7070D6B4F6E181C2 (IA6BBDC90BCC6EF2E35BFA8D709343BF3 ),
.I38B1AC532E13E69B05492C67EC7070BB (I5631F39935597168A2C9D3656C66CB5C ), .I705C64753A50CDA034B5ACB332D71768 (I0E620501249C5CFBF447631D04D33715 ),
.I233E0C0C8E5150F0CD8258F276D93942 ( ), .I102322A55721851004CB8E1F6AB50BDE (I25891FD4BF8EA7F9051CE324A21ED31E ),
.IBE0D6810EBD63B5C428623C578CF6D3A (I366EB0B781FD462E1BDC374519E76C20 ), .I115E90220158F08B0465E99D7F2561D3 ( )
); pmi_ram_dp # ( .pmi_wr_addr_depth (IB71844FFA3AB85FEF45EAB4D35395752 ), .pmi_wr_addr_width (I36A1B4EB5B5564A6ED7EA4D42856EFB4 ),
.pmi_wr_data_width (IF35F7B506981B2912E2486B227CB8871 ), .pmi_rd_addr_depth (IB71844FFA3AB85FEF45EAB4D35395752 ),
.pmi_rd_addr_width (I36A1B4EB5B5564A6ED7EA4D42856EFB4 ), .pmi_rd_data_width (IF35F7B506981B2912E2486B227CB8871 ),
.pmi_regmode ("reg"), .pmi_family (I66C185998F46A7148163982E39BCD296 ), .module_type ("pmi_ram_dp") )  I32900CECD80193336B4F376406D5DFF6
( .Data (IFD939E5BC1AA3DCE57CCDC18CA4F72A8 ), .RdAddress (IC2A6ECC367E2C82B97E73A57A8A79E1A ), .RdClockEn (1'b1),
.RdClock (ICCFB0F435B37370076102F325BC08D20 ), .Reset (I4AE98FF3DA4D5A5EE68F8A14D9D781F4 ), .WE (I25891FD4BF8EA7F9051CE324A21ED31E ),
.WrAddress (I5631F39935597168A2C9D3656C66CB5C ), .WrClockEn (1'b1), .WrClock (ICCFB0F435B37370076102F325BC08D20 ),
.Q (I2CA1A324143051A0AFDEFB54659C657C ) ); I4A464F8B941F768B40777E11E08CF0DE # ( .I7292F55C07BFD7FB8A60D29FFC186275
(I7292F55C07BFD7FB8A60D29FFC186275 ), .IDB9D60794264C5F8E5363941194A797B (IDB9D60794264C5F8E5363941194A797B ), .ID7C7F9F2E39BEBEE2ACFA8040034E48D
(ID7C7F9F2E39BEBEE2ACFA8040034E48D ) )  IC04A0BD824E0F4065A39094302E4599A ( .I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ),
.ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .IAB4F3026BD4F2760154E70C5BC0FE751 (I0E620501249C5CFBF447631D04D33715 ),
.ID8E639B3434FEAB4D1CA5AF230310D49 (I081545483B2E87A5F84E4E80F8AD87A7 ), .IC43B0BCCD0A723BBF62FF7B9D230C3F8 (I60B15FF62AA99717C8B7DA7D6912D281 ),
.I122CA37F449B813A5F0CAF8BC20EE9EA (I366EB0B781FD462E1BDC374519E76C20 ), .IFD5EF944B5EFFB20EE3422B3D79A2BF4 (ICB86B570A185B89048AE76A09444BA41 ),
.IB7C0B3EE4A87531F21610094A69146A7 (IE43DA634E45C0D88369455568042AF37 ), .IF87783FDF111A8E49EAC36F1DDFCBA80 (IF87783FDF111A8E49EAC36F1DDFCBA80 ),
.IF9D5978BE23690B1D4D13EF2AD676C6F (IF9D5978BE23690B1D4D13EF2AD676C6F ), .IDC6EA54AB52AEAD439CEF7521615AE1B (IDC6EA54AB52AEAD439CEF7521615AE1B ),
.I6ED49B5BED4BA586759FFDCC7B3B7FF8 (I6ED49B5BED4BA586759FFDCC7B3B7FF8 ), .I8E2F7CF6E50B95A483351A1836EB23AC (I8E2F7CF6E50B95A483351A1836EB23AC ),
.I506D2FCB600E0189274870B654E65B64 (I506D2FCB600E0189274870B654E65B64 ), .I141300E29D7EF4A0D8B71CB7469A7B90 (I141300E29D7EF4A0D8B71CB7469A7B90 ),
.I9AF8DD3F367CE82DF45437DB546EAAD3 (I9AF8DD3F367CE82DF45437DB546EAAD3 ), .I42D281FF99DC79A9AD9E7DF0AEB073A7 (I42D281FF99DC79A9AD9E7DF0AEB073A7 ),
.I3068B33EE97A971AE7F0CF17705AA6DC (I3068B33EE97A971AE7F0CF17705AA6DC ), .IFCBA19703D55B4610B3F4174C5B8833A (IFCBA19703D55B4610B3F4174C5B8833A ),
.IC3CC91D317012C130AC9E2A126F71C64 (IC3CC91D317012C130AC9E2A126F71C64 ), .ID8C32104758E11D83079BB9AEE0C35DB (I76EFAFF6D4391A79F5CD2CA7904431E8 ),
.IC91681A00788ED1B6C6956634033ED38 (IAFB0D72A35BE81312B83F6EC64D8ECF4 ), .I7114A89BF31DB18ED21FF0608A9BF50A (I9AC67CC0D048C17AC2F808C22F4DEE6F ),
.IB2B35E1DF060E7BC2B7E414954F6FA34 (IFD939E5BC1AA3DCE57CCDC18CA4F72A8 ), .I561BE0F01153FC1AADDEB08B34B545B6 (I6EFB980269078EDFE25D9139188C0357 ),
.IB86AF6EBEEA3CE1BF22AE1AF7CC8481F (ID6BA376F6FDCA561D55334C951D81896 ), .I94E3D00BBC13BF182097A25D63288C2C (I1261C037D95D7AC9FB55409369EA711E ),
.I8B25F4450817FC10E1E3DC6B500C9F5A (IAB4361F44053B3532F19F9BCB33E265F ), .I26C902CE18647F75561AD003E260B048 (I51F8ACA4F6E2B0688214E337318D090C ),
.IA5CEBFC654EDCA4107594F388D5BC88A (IAC7F9C0E3110EC41B40E14F4AFDB4D41 ), .I27627079DD78A85D26D85DC0C53D835F (I3645064ACD6F902F18DE49FBB6F7350B ),
.I0205131FB84BB0F9F8AD5CC00E5E861D (I64F37E01600233FCC804B26C0900CDE5 ), .IDA581E8478C8224118EF4E6B8EE8DDFE (ICA81D2D21EB4C7C4D7C6096277C9D15A ),
.IA36C0DD0DE88B03FA61EF35103D22DF0 (I200E0F93328C05371EF92973FC08E636 ) ); I2AA06444A0CB39074E17E74C913F2C98 #(
.I7292F55C07BFD7FB8A60D29FFC186275 (I7292F55C07BFD7FB8A60D29FFC186275 ), .I61D0345D311EC6FFC08DDDECE5F6127A (IB71844FFA3AB85FEF45EAB4D35395752 )
) ID1457574CA084B158A41B84E87670987 ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .IC79EC9A9F373F4B71374BDF6EDD31DE6 (1'b0), .ICFCA96AB1A120108CD0A9879E0F76EA8
(I2CA1A324143051A0AFDEFB54659C657C ), .ID8853B025150C80EE45BBA98E5BEA3A8 (I76EFAFF6D4391A79F5CD2CA7904431E8 ), .IF74C86FAF44E1757FDA146FCB1E10641
(I9AC67CC0D048C17AC2F808C22F4DEE6F ), .IA35D59E2E0D340C8C3D5ADB905E70579 (IA6BBDC90BCC6EF2E35BFA8D709343BF3 ), .I125028C7446331521D0434C10E8B0007
(I081545483B2E87A5F84E4E80F8AD87A7 ), .I0D04F33C419DDB2EC0886F4409AB9A96 (IE664D85E83E89DA36250C2ADD2CC9541 ), .I585F74DE05DD9C1C7070D6B4F6E181C2
(IE43DA634E45C0D88369455568042AF37 ) ); endmodule
 module IC067A254D727EC6E4653DEA8E2C9ED79 # (parameter I7292F55C07BFD7FB8A60D29FFC186275 = 32, parameter I7AEDD61970E812FD2535263A0E289FED
= 1, parameter I8B77F944A8EB2E113F742B8CB46E022C = 512, parameter I5A1D0B7A4A119DC7A35D6729D171C67D = 512, parameter
ICFA9960F43620DB191960C5C79DBFAE6 = 512, parameter IFB129920FFBFCFD17ADB3180F882E8E1 = 48 ) ( input wire ICCFB0F435B37370076102F325BC08D20 ,
input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire [7:0] IC680604FB338D55088F12313CDF2B03E , input wire [7:0]
IF17B1273FDE2637DBFCD3D142F80E5D5 , input wire [4:0] I44E00CA48D123AE945CB7C612A95BFE6 , input wire [2:0] I6D124B4E6D5F74B43E94949DE1CF46AA ,
input wire [2:0] I5C266315A3CF63C3FE988BB363C59AA1 , input wire [$clog2(I8B77F944A8EB2E113F742B8CB46E022C + 1) -
1:0] I8CE6978D396548B0C476A4C080ABF3CE , input wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] I879F5E0177BDD71945AEE80557DB31DC ,
input wire I3A0EE7E545E3C70F94B216D1405744A1 , input wire [$clog2(I5A1D0B7A4A119DC7A35D6729D171C67D + 1) - 1:0]
I7B58D405D154321FAF23051CBA4F0967 , input wire I2FBCFC2E8A11BEE681E33A995F23A9F7 , input wire I3EEFAC16E2400143CD0547F03531871C ,
input wire I7AC0939DFAAFF38545186E63551C4452 , input wire I9B878433B3D496FFA97B2BB22F930D6C , input wire [I7292F55C07BFD7FB8A60D29FFC186275
- 1:0] I886DDC9EB90AFC1350E4197DB0F9F21D , input wire IF63E3E7F031C0543230C8FA94864719C , input wire I081430FC44E0C370F3B3B4FAFFC51A69 ,
input wire [$clog2(ICFA9960F43620DB191960C5C79DBFAE6 + 1) - 1:0] I3FF97406B3ED373B267711109A980AF9 , input wire
I238A13C6F03704581F9A0A170F852FB4 , input wire I24C403550AE065D7D1B7266142886226 , input wire [IFB129920FFBFCFD17ADB3180F882E8E1
- 1:0] IDC6EA54AB52AEAD439CEF7521615AE1B , input wire [1:0] IC93EB5988EC451F72626A919FE396C61 , input wire [2:0]
I6ED49B5BED4BA586759FFDCC7B3B7FF8 , input wire [7:0] I8E2F7CF6E50B95A483351A1836EB23AC , input wire [I7292F55C07BFD7FB8A60D29FFC186275
- 1:0] I506D2FCB600E0189274870B654E65B64 , input wire [(I7292F55C07BFD7FB8A60D29FFC186275 / 8) - 1:0] I1304D1B0EBC59FFD53EF6CD7A8537E4D ,
input wire I141300E29D7EF4A0D8B71CB7469A7B90 , input wire IC3CC91D317012C130AC9E2A126F71C64 , output wire [7:0]
I7244B3A041E4EF91034ED304D36B4585 , output wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] I37622C557C24CD88B10BAD5A6CB7A4F4 ,
output wire I1E2C39A87E460C8AD520B4134F92292F , output wire I406DAF97F28CB5044A320565BE60692E , output wire ID24A83D781EA7F2CED8B0B12FADF20A5 ,
output wire IBADF395C0E67BC1FE7946C3D677241C4 , output wire IFB8B86C094497D5E859750490AB93CB4 , output wire IC3E8DB22A270F4E2527F04E7E81EFA46 ,
output wire IAEC671D12B80E2CC6E3D591A98E27230 , output wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] IA449B4CEADDC750F5446E3B900C14AA4 ,
output wire IFA413F55A4E38AA4A08DC60DCCB7553D , output wire I80F26623B387879BCA3F00C252D0129E , output wire [I7292F55C07BFD7FB8A60D29FFC186275
- 1:0] IFC7E490A5AF630CDD63895FB063ABE29 , output wire IEBE9989B3828CC1007CD10E6FBB2E76C , output wire I270ED686C2EF2C1C8B5B55EC4A5AAE84 ,
output wire IDA581E8478C8224118EF4E6B8EE8DDFE , output wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] I197028CF3B48BF15266050E66E13618E
);  `include "pcisig_constants.v" 
`include "wishbone_utils.v"
 localparam I2CDCB953A72C9DDCD6EF4FBE3D0BE88E = $clog2(I8B77F944A8EB2E113F742B8CB46E022C + 1); localparam IAB725F25E18FAFD445CA3B0B334590BE
= $clog2(I8B77F944A8EB2E113F742B8CB46E022C + 1); localparam I5D4944FED2815A3ECA7288050D4CB542 = IFB129920FFBFCFD17ADB3180F882E8E1
- 12; localparam IA056974EFE34F4C8FA362A54BD5FADF2 = 3; localparam IA948DD480C35DCCB0487F4F8B67FF99E = IFB129920FFBFCFD17ADB3180F882E8E1
- 1; localparam I1FC9733A3AF352A0F0C16A9487D3136E = 64 - IFB129920FFBFCFD17ADB3180F882E8E1 ; localparam [10:0] IF396FE43F94B3686844C6D5D6B5DB39C
= 11'b11111100000; localparam [10:0] IEBB19F00FE29431904C9AD7AC59816C6 = 11'b00000100000;  localparam IF8755D15B189AE86A6FDC2D1268FCDC9
= 6; localparam I24D2BA366F4F0CB889C7CBF7DBB156B6 = 6'b000000, I338F33967149E9BE8565EBC5277253E2 = 6'b000001, IE00763002B8F98799C282F18528369B1
= 6'b010000, I336B0D97AA4E31C1018007C9D81EE360 = 6'b010001, I5E31CC72F42872CA7609E04E3972135F = 6'b010010, I4E897662DE7109083665F92832975A0D
= 6'b010011, IFC5E1B899DC7A52E3A6263C63F5D7FBC = 6'b010100, I0AF4505AEE10B606D99FEB47577B3005 = 6'b010101, I1E0072D145F0522862103977C7AD48B5
= 6'b010110, ID89F181E16F6B4961901DD6C00C4FC50 = 6'b010111, I14E4373552472C84EAF0F2078975D1B7 = 6'b011000, IF5A542CAEF91CCA7EF42D20355D8815F
= 6'b100000, I1D81EEBBCFB3FB87EF20A35DFA862E9E = 6'b100001, I962095C6760357B792D0CD1278B21AF5 = 6'b100010, I9C2516A2CE92B199562345D5833785B3
= 6'b100011, I8A8F7A096F2E5012EDBEBDDEB9EEE34E = 6'b100100, IC6B19C3976DC11C4C29F6DFCC51BB3CF = 6'b100101, I11ABAF7FCD68013E37F52A8A41493B59
= 6'b100110, I3FC158820A9D44CAF3F67A39EBCD3D14 = 6'b100111, IEA810C9EE9AC978D2DFB6A0C31191743 = 6'b101000;  reg
[9:0] I0CE969690E7FBD3AD68AAD352783F26A ; reg [3:0] I11FD35FED78BCB8861FACB9A1E3A4C35 ; reg [3:0] IC52F3B77F7E45A74323561D6A6F6028A ;
reg [7:0] IBA8C2E9643A807EAD24886E1C89ED4E1 ; reg IF4B2F356412545C21578876129150C2F ; reg [10:0] ID5D5AB03A95A35F722F49CD4B0E185F1 ;
reg [2:0] I2792804BC0B8F3DDCC1D08D4DE2F25DA ; reg [2:0] IE763761FF58557F78DA03BEF9DCF712E ; reg [10:0] I96151A81C6E1327A706028BA81B3E8AE ;
reg [7:0] I4C387EC384562841515F49E7547AFA1E ; reg I2B169A80A1410659B701DC07563639A3 ; reg IFFBEF8AE96EE878792DDB3FCC731CB4B ;
reg I1E515C54DF69EFC5334ACB78A7F46488 ; reg I0DE270F6B1F18A35E6835C0695437A55 ; reg IBCBE72A344F91A6C63C524CD8C9FFBAC ;
reg [10:0] I0B6ECB7D58876821FA73D9499B8DE015 ; reg I6425A964B876A53D38FE4C91B5A930BF ; reg [31:0] I81CA76177EADF878D9C5F8B834BC9401 ;
reg I62FE0E7DC25E3D62EEE0FBBDF869D2E8 ; reg IF9EE6A022EB9CA07758C3F88273952CB ; reg [10:0] IEB5C97BD73E9C46378468349D65DB2D9 ;
reg [9:0] I494F8E6C428E0D5AB7D0135AD31F3C46 ; reg [10:0] I3EC90F87E70407C2A46DA25A8CA9065B ; reg I87570FA9CFC0EF2B57A30C0D3942AD58 ;
reg IF3EB173FF5CCD07FA7EB0E8A13FE3FE3 ; reg I9DF7D0AF404EC4CE8D1499B20F238C23 ; reg [31:0] I77B1E95A01761A9A5D153F6B403BCE8E ;
reg IFFD521EABA6F14D35240B97DD5930909 ; reg I4146C7DC49C187159B0A3C9D44515C29 ; reg IEE09BFC6815DBA057FA2D268AD02EFDA ;
reg IE44E1C3E3A8A49BF1C8E3C7ADFBE8CD5 ; reg I670A86ADD4DA92DA04F0354154D50812 ; reg IA42493546F7BB75836172B5E62E7CDF2 ;
reg I8D181359467F27637239CDAEE8A2F45A ; reg IF58956C1F9E72353D1F5C742AE29FB85 ; reg IA30591CFD911D315F76A63BA264689D4 ;
reg I5A09FE74EFC8C7CD279F9D32F0E4BF2A ; reg [9:0] ICED1EF5C0E5400F7869E1C674AE21DA6 ; reg [7:0] ID564A30F71C7C1B827BA57264E89B21D ;
reg [31:0] I44109A75F9883AA09218902DA5B2CBB3 ; reg [31:0] I074FD9C5AE408613B3750B75A6125486 ; reg [2:0] I5FC6334EB24FE23F5733F744B8E73624 ;
reg [I5D4944FED2815A3ECA7288050D4CB542 - 1:0] IE48F23B4AE45A1E423AC11ED564DE4D8 ; reg [9:0] IABB783BAEC6EC4928216CD800CAC26FC ;
reg [9:0] I83C959FA1B0FD40F9B8261F8DA6D2791 ; reg I21AD57B50E491E60E17CBE10D72C4241 ; reg I36FECBB048E15937DC767259CBABEDCB ;
reg [IF8755D15B189AE86A6FDC2D1268FCDC9 - 1:0] I706E9793A36552E97EF7B1CF0F6162D7 ; reg [IF8755D15B189AE86A6FDC2D1268FCDC9
- 1:0] I1915785CFF3E5F70FE78AAE0F38632BE ; wire I6D75D178107F34EC234BF34C357BEAE3 ; wire I3DA025A250DA8401A3758BF5C2D7CF37 ;
wire IA28DF69CCCF33F049890BA79F1203E18 ; wire I61BE5C1B2846DC2A3D30184D92B188B0 ; wire I39897CE0B696B5ACFB39C404E7230CD4 ;
wire I2D3F6195192E51E825219F43C080A709 ; wire IFC805C60848CB0108E26B68757DC3B62 ; wire IEA2F6215D00C222A05E71C8508532AB0 ;
wire IB5358AE45A21CC9091163666F5E272C8 ;  assign I7244B3A041E4EF91034ED304D36B4585 = I4C387EC384562841515F49E7547AFA1E ;
assign I37622C557C24CD88B10BAD5A6CB7A4F4 = I44109A75F9883AA09218902DA5B2CBB3 ; assign I1E2C39A87E460C8AD520B4134F92292F
= IBCBE72A344F91A6C63C524CD8C9FFBAC ; assign I406DAF97F28CB5044A320565BE60692E = I3DA025A250DA8401A3758BF5C2D7CF37 ;
assign ID24A83D781EA7F2CED8B0B12FADF20A5 = I6425A964B876A53D38FE4C91B5A930BF ; assign IBADF395C0E67BC1FE7946C3D677241C4
= I9DF7D0AF404EC4CE8D1499B20F238C23 | I39897CE0B696B5ACFB39C404E7230CD4 ; assign IC3E8DB22A270F4E2527F04E7E81EFA46
= IFFD521EABA6F14D35240B97DD5930909 ; assign IAEC671D12B80E2CC6E3D591A98E27230 = I4146C7DC49C187159B0A3C9D44515C29 ;
assign IA449B4CEADDC750F5446E3B900C14AA4 = I77B1E95A01761A9A5D153F6B403BCE8E ; assign IFA413F55A4E38AA4A08DC60DCCB7553D
= IEE09BFC6815DBA057FA2D268AD02EFDA ; assign I80F26623B387879BCA3F00C252D0129E = I670A86ADD4DA92DA04F0354154D50812
| I62FE0E7DC25E3D62EEE0FBBDF869D2E8 ; assign IFC7E490A5AF630CDD63895FB063ABE29 = (I62FE0E7DC25E3D62EEE0FBBDF869D2E8 )
? I81CA76177EADF878D9C5F8B834BC9401 : I77B1E95A01761A9A5D153F6B403BCE8E ; assign IEBE9989B3828CC1007CD10E6FBB2E76C
= IA42493546F7BB75836172B5E62E7CDF2 ; assign I270ED686C2EF2C1C8B5B55EC4A5AAE84 = I8D181359467F27637239CDAEE8A2F45A ;
assign IFB8B86C094497D5E859750490AB93CB4 = 1'b0; assign IDA581E8478C8224118EF4E6B8EE8DDFE = I2D3F6195192E51E825219F43C080A709 ;
assign I197028CF3B48BF15266050E66E13618E = I074FD9C5AE408613B3750B75A6125486 ;  assign I6D75D178107F34EC234BF34C357BEAE3
= IFFBEF8AE96EE878792DDB3FCC731CB4B | I1E515C54DF69EFC5334ACB78A7F46488 ; assign I3DA025A250DA8401A3758BF5C2D7CF37
= (|I0B6ECB7D58876821FA73D9499B8DE015 ) & IE44E1C3E3A8A49BF1C8E3C7ADFBE8CD5 ; assign IA28DF69CCCF33F049890BA79F1203E18
= (I706E9793A36552E97EF7B1CF0F6162D7 == IEA810C9EE9AC978D2DFB6A0C31191743 ) ? IF9EE6A022EB9CA07758C3F88273952CB
: 1'b0; assign I61BE5C1B2846DC2A3D30184D92B188B0 = ~I83C959FA1B0FD40F9B8261F8DA6D2791 [0]; assign I39897CE0B696B5ACFB39C404E7230CD4
= (I706E9793A36552E97EF7B1CF0F6162D7 == I14E4373552472C84EAF0F2078975D1B7 ) ? ~IF63E3E7F031C0543230C8FA94864719C
: 1'b0; assign I2D3F6195192E51E825219F43C080A709 = IF58956C1F9E72353D1F5C742AE29FB85 | I5A09FE74EFC8C7CD279F9D32F0E4BF2A ;
assign IFC805C60848CB0108E26B68757DC3B62 = (I6ED49B5BED4BA586759FFDCC7B3B7FF8 == IEE94C2462F89091D3C62992327532D1E )
? IB5358AE45A21CC9091163666F5E272C8 : 1'b0; assign IEA2F6215D00C222A05E71C8508532AB0 = (I6ED49B5BED4BA586759FFDCC7B3B7FF8
== IEE94C2462F89091D3C62992327532D1E ) ? 1'b1 : 1'b0; assign IB5358AE45A21CC9091163666F5E272C8 = I2D3F6195192E51E825219F43C080A709
& I141300E29D7EF4A0D8B71CB7469A7B90 & (|I8E2F7CF6E50B95A483351A1836EB23AC );  always @(*) begin I1915785CFF3E5F70FE78AAE0F38632BE
= I706E9793A36552E97EF7B1CF0F6162D7 ; case (I706E9793A36552E97EF7B1CF0F6162D7 ) I24D2BA366F4F0CB889C7CBF7DBB156B6
: begin if (I8E2F7CF6E50B95A483351A1836EB23AC & IBA8C2E9643A807EAD24886E1C89ED4E1 ) I1915785CFF3E5F70FE78AAE0F38632BE
= I338F33967149E9BE8565EBC5277253E2 ; end I338F33967149E9BE8565EBC5277253E2 : begin if (I36FECBB048E15937DC767259CBABEDCB )
I1915785CFF3E5F70FE78AAE0F38632BE = IF5A542CAEF91CCA7EF42D20355D8815F ; else if (I2B169A80A1410659B701DC07563639A3 )
I1915785CFF3E5F70FE78AAE0F38632BE = IE00763002B8F98799C282F18528369B1 ; end IE00763002B8F98799C282F18528369B1 :
begin I1915785CFF3E5F70FE78AAE0F38632BE = I336B0D97AA4E31C1018007C9D81EE360 ; end I336B0D97AA4E31C1018007C9D81EE360
: begin I1915785CFF3E5F70FE78AAE0F38632BE = I5E31CC72F42872CA7609E04E3972135F ; end I5E31CC72F42872CA7609E04E3972135F
: begin I1915785CFF3E5F70FE78AAE0F38632BE = I4E897662DE7109083665F92832975A0D ; end I4E897662DE7109083665F92832975A0D
: begin I1915785CFF3E5F70FE78AAE0F38632BE = IFC5E1B899DC7A52E3A6263C63F5D7FBC ; end IFC5E1B899DC7A52E3A6263C63F5D7FBC
: begin if (IF4B2F356412545C21578876129150C2F ) I1915785CFF3E5F70FE78AAE0F38632BE = I0AF4505AEE10B606D99FEB47577B3005 ;
else I1915785CFF3E5F70FE78AAE0F38632BE = I1E0072D145F0522862103977C7AD48B5 ; end I0AF4505AEE10B606D99FEB47577B3005
: begin I1915785CFF3E5F70FE78AAE0F38632BE = I1E0072D145F0522862103977C7AD48B5 ; end I1E0072D145F0522862103977C7AD48B5
: begin if (I238A13C6F03704581F9A0A170F852FB4 ) I1915785CFF3E5F70FE78AAE0F38632BE = ID89F181E16F6B4961901DD6C00C4FC50 ;
end ID89F181E16F6B4961901DD6C00C4FC50 : begin if (~(|I3EC90F87E70407C2A46DA25A8CA9065B ) & IF63E3E7F031C0543230C8FA94864719C
& ~(|IEB5C97BD73E9C46378468349D65DB2D9 )) I1915785CFF3E5F70FE78AAE0F38632BE = I24D2BA366F4F0CB889C7CBF7DBB156B6 ;
else if (IFC805C60848CB0108E26B68757DC3B62 ) I1915785CFF3E5F70FE78AAE0F38632BE = I14E4373552472C84EAF0F2078975D1B7 ;
end I14E4373552472C84EAF0F2078975D1B7 : begin if (~(|I3EC90F87E70407C2A46DA25A8CA9065B ) & IF63E3E7F031C0543230C8FA94864719C
& ~I7AC0939DFAAFF38545186E63551C4452 & ~IF3EB173FF5CCD07FA7EB0E8A13FE3FE3 ) I1915785CFF3E5F70FE78AAE0F38632BE =
I24D2BA366F4F0CB889C7CBF7DBB156B6 ; end IF5A542CAEF91CCA7EF42D20355D8815F : begin if (IFC805C60848CB0108E26B68757DC3B62
| I6D75D178107F34EC234BF34C357BEAE3 ) if (IE44E1C3E3A8A49BF1C8E3C7ADFBE8CD5 & ~(|I0B6ECB7D58876821FA73D9499B8DE015 ))
I1915785CFF3E5F70FE78AAE0F38632BE = I962095C6760357B792D0CD1278B21AF5 ; else I1915785CFF3E5F70FE78AAE0F38632BE =
I1D81EEBBCFB3FB87EF20A35DFA862E9E ; end I1D81EEBBCFB3FB87EF20A35DFA862E9E : begin if (IE44E1C3E3A8A49BF1C8E3C7ADFBE8CD5
& ~(|I0B6ECB7D58876821FA73D9499B8DE015 )) I1915785CFF3E5F70FE78AAE0F38632BE = I962095C6760357B792D0CD1278B21AF5 ;
end I962095C6760357B792D0CD1278B21AF5 : begin I1915785CFF3E5F70FE78AAE0F38632BE = I9C2516A2CE92B199562345D5833785B3 ;
end I9C2516A2CE92B199562345D5833785B3 : begin I1915785CFF3E5F70FE78AAE0F38632BE = I8A8F7A096F2E5012EDBEBDDEB9EEE34E ;
end I8A8F7A096F2E5012EDBEBDDEB9EEE34E : begin if (IF4B2F356412545C21578876129150C2F ) I1915785CFF3E5F70FE78AAE0F38632BE
= IC6B19C3976DC11C4C29F6DFCC51BB3CF ; else I1915785CFF3E5F70FE78AAE0F38632BE = I11ABAF7FCD68013E37F52A8A41493B59 ;
end IC6B19C3976DC11C4C29F6DFCC51BB3CF : begin I1915785CFF3E5F70FE78AAE0F38632BE = I11ABAF7FCD68013E37F52A8A41493B59 ;
end    I11ABAF7FCD68013E37F52A8A41493B59 : begin if (I21AD57B50E491E60E17CBE10D72C4241 ) I1915785CFF3E5F70FE78AAE0F38632BE
= I3FC158820A9D44CAF3F67A39EBCD3D14 ; else I1915785CFF3E5F70FE78AAE0F38632BE = IF5A542CAEF91CCA7EF42D20355D8815F ;
end I3FC158820A9D44CAF3F67A39EBCD3D14 : begin if (~(|I0B6ECB7D58876821FA73D9499B8DE015 ) & ~I2FBCFC2E8A11BEE681E33A995F23A9F7 )
I1915785CFF3E5F70FE78AAE0F38632BE = IEA810C9EE9AC978D2DFB6A0C31191743 ; end IEA810C9EE9AC978D2DFB6A0C31191743 :
begin if (I24C403550AE065D7D1B7266142886226 ) I1915785CFF3E5F70FE78AAE0F38632BE = I24D2BA366F4F0CB889C7CBF7DBB156B6 ;
end default : begin end endcase end  always @(posedge ICCFB0F435B37370076102F325BC08D20 or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 )
begin if (~I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin I0CE969690E7FBD3AD68AAD352783F26A <= 10'b0; I11FD35FED78BCB8861FACB9A1E3A4C35
<= 4'b0; IC52F3B77F7E45A74323561D6A6F6028A <= 4'b0; IBA8C2E9643A807EAD24886E1C89ED4E1 <= 8'b0; IF4B2F356412545C21578876129150C2F
<= 1'b0; ID5D5AB03A95A35F722F49CD4B0E185F1 <= 11'b0; I2792804BC0B8F3DDCC1D08D4DE2F25DA <= 3'b0; IE763761FF58557F78DA03BEF9DCF712E
<= 3'b0; I96151A81C6E1327A706028BA81B3E8AE <= 11'b0; I4C387EC384562841515F49E7547AFA1E <= 8'b0; I2B169A80A1410659B701DC07563639A3
<= 1'b0; IFFBEF8AE96EE878792DDB3FCC731CB4B <= 1'b0; I1E515C54DF69EFC5334ACB78A7F46488 <= 1'b0; IBCBE72A344F91A6C63C524CD8C9FFBAC
<= 1'b0; I0B6ECB7D58876821FA73D9499B8DE015 <= 11'b0; I6425A964B876A53D38FE4C91B5A930BF <= 1'b0; I0DE270F6B1F18A35E6835C0695437A55
<= 1'b0; I81CA76177EADF878D9C5F8B834BC9401 <= 32'b0; I62FE0E7DC25E3D62EEE0FBBDF869D2E8 <= 1'b0; IF9EE6A022EB9CA07758C3F88273952CB
<= 1'b0; IFFD521EABA6F14D35240B97DD5930909 <= 1'b0; I4146C7DC49C187159B0A3C9D44515C29 <= 1'b0; IEE09BFC6815DBA057FA2D268AD02EFDA
<= 1'b0; IE44E1C3E3A8A49BF1C8E3C7ADFBE8CD5 <= 1'b0; I670A86ADD4DA92DA04F0354154D50812 <= 1'b0; IEB5C97BD73E9C46378468349D65DB2D9
<= 11'b0; I494F8E6C428E0D5AB7D0135AD31F3C46 <= 10'b0; I3EC90F87E70407C2A46DA25A8CA9065B <= 11'b0; IF3EB173FF5CCD07FA7EB0E8A13FE3FE3
<= 1'b0; I9DF7D0AF404EC4CE8D1499B20F238C23 <= 1'b0; I77B1E95A01761A9A5D153F6B403BCE8E <= 32'b0; IA42493546F7BB75836172B5E62E7CDF2
<= 1'b0; I8D181359467F27637239CDAEE8A2F45A <= 1'b0; IF58956C1F9E72353D1F5C742AE29FB85 <= 1'b0; IA30591CFD911D315F76A63BA264689D4
<= 1'b0; I5A09FE74EFC8C7CD279F9D32F0E4BF2A <= 1'b0; ICED1EF5C0E5400F7869E1C674AE21DA6 <= 10'b0; ID564A30F71C7C1B827BA57264E89B21D
<= 8'b0; I44109A75F9883AA09218902DA5B2CBB3 <= 32'b0; I074FD9C5AE408613B3750B75A6125486 <= 32'b0; I5FC6334EB24FE23F5733F744B8E73624
<= 3'b0; IE48F23B4AE45A1E423AC11ED564DE4D8 <= {I5D4944FED2815A3ECA7288050D4CB542 {1'b0}}; IABB783BAEC6EC4928216CD800CAC26FC
<= 10'b0; I83C959FA1B0FD40F9B8261F8DA6D2791 <= 10'b0; I21AD57B50E491E60E17CBE10D72C4241 <= 1'b0; I36FECBB048E15937DC767259CBABEDCB
<= 1'b0; I706E9793A36552E97EF7B1CF0F6162D7 <= I24D2BA366F4F0CB889C7CBF7DBB156B6 ; end else begin I0CE969690E7FBD3AD68AAD352783F26A
<= IF396FE43F94B3686844C6D5D6B5DB39C << IE763761FF58557F78DA03BEF9DCF712E ; IBA8C2E9643A807EAD24886E1C89ED4E1 <=
IC680604FB338D55088F12313CDF2B03E ; IE763761FF58557F78DA03BEF9DCF712E <= I5C266315A3CF63C3FE988BB363C59AA1 ; I96151A81C6E1327A706028BA81B3E8AE
<= IEBB19F00FE29431904C9AD7AC59816C6 << IE763761FF58557F78DA03BEF9DCF712E ; I4C387EC384562841515F49E7547AFA1E <=
I8E2F7CF6E50B95A483351A1836EB23AC ; IBCBE72A344F91A6C63C524CD8C9FFBAC <= 1'b0; I6425A964B876A53D38FE4C91B5A930BF
<= (I706E9793A36552E97EF7B1CF0F6162D7 == IF5A542CAEF91CCA7EF42D20355D8815F ) ? IB5358AE45A21CC9091163666F5E272C8
: 1'b0; I81CA76177EADF878D9C5F8B834BC9401 <= {I879F5E0177BDD71945AEE80557DB31DC [7:0], I879F5E0177BDD71945AEE80557DB31DC [15:8],
I879F5E0177BDD71945AEE80557DB31DC [23:16], I879F5E0177BDD71945AEE80557DB31DC [31:24]}; I62FE0E7DC25E3D62EEE0FBBDF869D2E8
<= I2FBCFC2E8A11BEE681E33A995F23A9F7 | IA28DF69CCCF33F049890BA79F1203E18 ; I494F8E6C428E0D5AB7D0135AD31F3C46 <=
I96151A81C6E1327A706028BA81B3E8AE [9:0] - (IABB783BAEC6EC4928216CD800CAC26FC & ~I0CE969690E7FBD3AD68AAD352783F26A [9:0]);
IF3EB173FF5CCD07FA7EB0E8A13FE3FE3 <= I7AC0939DFAAFF38545186E63551C4452 ; IFFD521EABA6F14D35240B97DD5930909 <= 1'b0;
I4146C7DC49C187159B0A3C9D44515C29 <= 1'b0; IEE09BFC6815DBA057FA2D268AD02EFDA <= (I7AEDD61970E812FD2535263A0E289FED
== 1) ? I3A0EE7E545E3C70F94B216D1405744A1 : ((IF9EE6A022EB9CA07758C3F88273952CB ) ? IA28DF69CCCF33F049890BA79F1203E18
: I3A0EE7E545E3C70F94B216D1405744A1 ); I670A86ADD4DA92DA04F0354154D50812 <= 1'b0; I2B169A80A1410659B701DC07563639A3
<= (I8CE6978D396548B0C476A4C080ABF3CE > 3) ? 1'b1 : 1'b0; I0DE270F6B1F18A35E6835C0695437A55 <= (I7B58D405D154321FAF23051CBA4F0967
> IA056974EFE34F4C8FA362A54BD5FADF2 ) ? 1'b1 : 1'b0; IE44E1C3E3A8A49BF1C8E3C7ADFBE8CD5 <= (I3FF97406B3ED373B267711109A980AF9
> 3) ? 1'b1 : 1'b0; I9DF7D0AF404EC4CE8D1499B20F238C23 <= ~I36FECBB048E15937DC767259CBABEDCB & ~(I9DF7D0AF404EC4CE8D1499B20F238C23
& I9B878433B3D496FFA97B2BB22F930D6C ) & ~I21AD57B50E491E60E17CBE10D72C4241 & ((~IF63E3E7F031C0543230C8FA94864719C
& ~IF58956C1F9E72353D1F5C742AE29FB85 ) | (~IF63E3E7F031C0543230C8FA94864719C & IB5358AE45A21CC9091163666F5E272C8
& ~IFC805C60848CB0108E26B68757DC3B62 )); I5A09FE74EFC8C7CD279F9D32F0E4BF2A <= 1'b0; I21AD57B50E491E60E17CBE10D72C4241
<= (I706E9793A36552E97EF7B1CF0F6162D7 == I338F33967149E9BE8565EBC5277253E2 ) ? 1'b0 : (I21AD57B50E491E60E17CBE10D72C4241
| IFC805C60848CB0108E26B68757DC3B62 ); I706E9793A36552E97EF7B1CF0F6162D7 <= I1915785CFF3E5F70FE78AAE0F38632BE ;
if (I7AC0939DFAAFF38545186E63551C4452 ) I3EC90F87E70407C2A46DA25A8CA9065B <= (I3EC90F87E70407C2A46DA25A8CA9065B
< I7AEDD61970E812FD2535263A0E289FED ) ? 0 : (I3EC90F87E70407C2A46DA25A8CA9065B - I7AEDD61970E812FD2535263A0E289FED );
if (|I0B6ECB7D58876821FA73D9499B8DE015 ) begin if (I3DA025A250DA8401A3758BF5C2D7CF37 ) I0B6ECB7D58876821FA73D9499B8DE015
<= I0B6ECB7D58876821FA73D9499B8DE015 - 1; end if (IFC805C60848CB0108E26B68757DC3B62 ) begin I074FD9C5AE408613B3750B75A6125486
<= 32'b0; IF58956C1F9E72353D1F5C742AE29FB85 <= 1'b0; end else begin IF58956C1F9E72353D1F5C742AE29FB85 <= (I081430FC44E0C370F3B3B4FAFFC51A69
& ~I21AD57B50E491E60E17CBE10D72C4241 & ~IA30591CFD911D315F76A63BA264689D4 ) | (IF58956C1F9E72353D1F5C742AE29FB85
& ~IB5358AE45A21CC9091163666F5E272C8 ); IA30591CFD911D315F76A63BA264689D4 <= IA30591CFD911D315F76A63BA264689D4 &
~I081430FC44E0C370F3B3B4FAFFC51A69 ; if (I081430FC44E0C370F3B3B4FAFFC51A69 ) I074FD9C5AE408613B3750B75A6125486 <=
I886DDC9EB90AFC1350E4197DB0F9F21D ; end  case (I706E9793A36552E97EF7B1CF0F6162D7 ) I5E31CC72F42872CA7609E04E3972135F
: begin IEB5C97BD73E9C46378468349D65DB2D9 <= {~(|I494F8E6C428E0D5AB7D0135AD31F3C46 ), I494F8E6C428E0D5AB7D0135AD31F3C46 };
end I14E4373552472C84EAF0F2078975D1B7 : begin IEB5C97BD73E9C46378468349D65DB2D9 <= 11'b0; end default : begin IEB5C97BD73E9C46378468349D65DB2D9
<= (IEB5C97BD73E9C46378468349D65DB2D9 && IB5358AE45A21CC9091163666F5E272C8 ) ? IEB5C97BD73E9C46378468349D65DB2D9
- 1 : IEB5C97BD73E9C46378468349D65DB2D9 ; end endcase  case (I706E9793A36552E97EF7B1CF0F6162D7 ) I24D2BA366F4F0CB889C7CBF7DBB156B6
: begin if (I8E2F7CF6E50B95A483351A1836EB23AC ) begin I11FD35FED78BCB8861FACB9A1E3A4C35 <= I1304D1B0EBC59FFD53EF6CD7A8537E4D ;
I2792804BC0B8F3DDCC1D08D4DE2F25DA <= I6D124B4E6D5F74B43E94949DE1CF46AA ; ID564A30F71C7C1B827BA57264E89B21D <= I8E2F7CF6E50B95A483351A1836EB23AC ;
I36FECBB048E15937DC767259CBABEDCB <= IC3CC91D317012C130AC9E2A126F71C64 ; end end I338F33967149E9BE8565EBC5277253E2
: begin IC52F3B77F7E45A74323561D6A6F6028A <= 4'b0; IFFBEF8AE96EE878792DDB3FCC731CB4B <= &IDC6EA54AB52AEAD439CEF7521615AE1B [11:2];
I1E515C54DF69EFC5334ACB78A7F46488 <= 1'b0; I5A09FE74EFC8C7CD279F9D32F0E4BF2A <= I0DE270F6B1F18A35E6835C0695437A55
& I36FECBB048E15937DC767259CBABEDCB ; ICED1EF5C0E5400F7869E1C674AE21DA6 <= 1; I21AD57B50E491E60E17CBE10D72C4241
<= 1'b0; {IE48F23B4AE45A1E423AC11ED564DE4D8 , IABB783BAEC6EC4928216CD800CAC26FC } <= IDC6EA54AB52AEAD439CEF7521615AE1B [IA948DD480C35DCCB0487F4F8B67FF99E :2];
I83C959FA1B0FD40F9B8261F8DA6D2791 <= IDC6EA54AB52AEAD439CEF7521615AE1B [11:2]; case (I2792804BC0B8F3DDCC1D08D4DE2F25DA )
1 : begin ID5D5AB03A95A35F722F49CD4B0E185F1 <= 11'd64; end 2 : begin ID5D5AB03A95A35F722F49CD4B0E185F1 <= 11'd128;
end 3 : begin ID5D5AB03A95A35F722F49CD4B0E185F1 <= 11'd256; end 4 : begin ID5D5AB03A95A35F722F49CD4B0E185F1 <= 11'd512;
end 5 : begin ID5D5AB03A95A35F722F49CD4B0E185F1 <= 11'd1024; end default : begin ID5D5AB03A95A35F722F49CD4B0E185F1
<= 11'd32; end endcase case (ID564A30F71C7C1B827BA57264E89B21D ) 8'h02 : begin I5FC6334EB24FE23F5733F744B8E73624
<= 3'h1; end 8'h04 : begin I5FC6334EB24FE23F5733F744B8E73624 <= 3'h2; end 8'h08 : begin I5FC6334EB24FE23F5733F744B8E73624
<= 3'h3; end 8'h10 : begin I5FC6334EB24FE23F5733F744B8E73624 <= 3'h4; end 8'h20 : begin I5FC6334EB24FE23F5733F744B8E73624
<= 3'h5; end 8'h40 : begin I5FC6334EB24FE23F5733F744B8E73624 <= 3'h6; end 8'h80 : begin I5FC6334EB24FE23F5733F744B8E73624
<= 3'h7; end default : begin I5FC6334EB24FE23F5733F744B8E73624 <= 3'h0; end endcase end IE00763002B8F98799C282F18528369B1
: begin I11FD35FED78BCB8861FACB9A1E3A4C35 <= {4{1'b1}}; IF4B2F356412545C21578876129150C2F <= |(IE48F23B4AE45A1E423AC11ED564DE4D8 [I5D4944FED2815A3ECA7288050D4CB542
- 1:20]); IA30591CFD911D315F76A63BA264689D4 <= (I7AEDD61970E812FD2535263A0E289FED > 1) ? I83C959FA1B0FD40F9B8261F8DA6D2791 [0]
: 1'b0; end I336B0D97AA4E31C1018007C9D81EE360 : begin I3EC90F87E70407C2A46DA25A8CA9065B [9:0] <= I494F8E6C428E0D5AB7D0135AD31F3C46 ;
I3EC90F87E70407C2A46DA25A8CA9065B [10] <= ~(|I494F8E6C428E0D5AB7D0135AD31F3C46 ); if (I494F8E6C428E0D5AB7D0135AD31F3C46
== 1) IC52F3B77F7E45A74323561D6A6F6028A <= {4{1'b0}}; else IC52F3B77F7E45A74323561D6A6F6028A <= {4{1'b1}}; end I5E31CC72F42872CA7609E04E3972135F
: begin I4146C7DC49C187159B0A3C9D44515C29 <= 1'b1; if (IF4B2F356412545C21578876129150C2F ) I77B1E95A01761A9A5D153F6B403BCE8E
<= {I877B2A234FC10EC8A4A2F0A90F6EAE6C , {14{1'b0}}, I494F8E6C428E0D5AB7D0135AD31F3C46 }; else I77B1E95A01761A9A5D153F6B403BCE8E
<= {I8F0EB88EC813DC0B3105F31BABD34B79 , {14{1'b0}}, I494F8E6C428E0D5AB7D0135AD31F3C46 }; end I4E897662DE7109083665F92832975A0D
: begin  I4146C7DC49C187159B0A3C9D44515C29 <= 1'b1; I77B1E95A01761A9A5D153F6B403BCE8E <= {IF17B1273FDE2637DBFCD3D142F80E5D5 ,
I44E00CA48D123AE945CB7C612A95BFE6 , I5FC6334EB24FE23F5733F744B8E73624 , {8{1'b0}}, IC52F3B77F7E45A74323561D6A6F6028A ,
I11FD35FED78BCB8861FACB9A1E3A4C35 }; end IFC5E1B899DC7A52E3A6263C63F5D7FBC : begin IFFD521EABA6F14D35240B97DD5930909
<= ~IF4B2F356412545C21578876129150C2F ; I4146C7DC49C187159B0A3C9D44515C29 <= 1'b1; if (IF4B2F356412545C21578876129150C2F )
I77B1E95A01761A9A5D153F6B403BCE8E <= {{I1FC9733A3AF352A0F0C16A9487D3136E {1'b0}}, IE48F23B4AE45A1E423AC11ED564DE4D8 [I5D4944FED2815A3ECA7288050D4CB542
- 1:20]}; else I77B1E95A01761A9A5D153F6B403BCE8E <= {IE48F23B4AE45A1E423AC11ED564DE4D8 [19:0], I83C959FA1B0FD40F9B8261F8DA6D2791 ,
{2{1'b0}}}; end I0AF4505AEE10B606D99FEB47577B3005 : begin IFFD521EABA6F14D35240B97DD5930909 <= 1'b1; I4146C7DC49C187159B0A3C9D44515C29
<= 1'b1; I77B1E95A01761A9A5D153F6B403BCE8E <= {IE48F23B4AE45A1E423AC11ED564DE4D8 [19:0], I83C959FA1B0FD40F9B8261F8DA6D2791 ,
{2{1'b0}}}; end I1E0072D145F0522862103977C7AD48B5 : begin IA42493546F7BB75836172B5E62E7CDF2 <= ~IA42493546F7BB75836172B5E62E7CDF2
| (IA42493546F7BB75836172B5E62E7CDF2 & ~I238A13C6F03704581F9A0A170F852FB4 ); end IF5A542CAEF91CCA7EF42D20355D8815F
: begin IF4B2F356412545C21578876129150C2F <= |(IE48F23B4AE45A1E423AC11ED564DE4D8 [I5D4944FED2815A3ECA7288050D4CB542
- 1:20]); if (I2D3F6195192E51E825219F43C080A709 & |I8E2F7CF6E50B95A483351A1836EB23AC & I141300E29D7EF4A0D8B71CB7469A7B90 )
begin IFFBEF8AE96EE878792DDB3FCC731CB4B <= &IABB783BAEC6EC4928216CD800CAC26FC [9:1]; I1E515C54DF69EFC5334ACB78A7F46488
<= (ICED1EF5C0E5400F7869E1C674AE21DA6 == (ID5D5AB03A95A35F722F49CD4B0E185F1 - 1)) ? 1'b1 : 1'b0; IBCBE72A344F91A6C63C524CD8C9FFBAC
<= I6D75D178107F34EC234BF34C357BEAE3 | IEA2F6215D00C222A05E71C8508532AB0 ; I5A09FE74EFC8C7CD279F9D32F0E4BF2A <=
(I0DE270F6B1F18A35E6835C0695437A55 ) ? (~ (IEA2F6215D00C222A05E71C8508532AB0 | I6D75D178107F34EC234BF34C357BEAE3 ))
: 1'b0; I44109A75F9883AA09218902DA5B2CBB3 <= I506D2FCB600E0189274870B654E65B64 ; IABB783BAEC6EC4928216CD800CAC26FC
<= IABB783BAEC6EC4928216CD800CAC26FC + 1; if (I6D75D178107F34EC234BF34C357BEAE3 | IEA2F6215D00C222A05E71C8508532AB0 )
IF9EE6A022EB9CA07758C3F88273952CB <= (I7AEDD61970E812FD2535263A0E289FED == 1) ? 1'b0 : (IF4B2F356412545C21578876129150C2F
? ICED1EF5C0E5400F7869E1C674AE21DA6 [0] : ~ICED1EF5C0E5400F7869E1C674AE21DA6 [0]); else ICED1EF5C0E5400F7869E1C674AE21DA6
<= ICED1EF5C0E5400F7869E1C674AE21DA6 + 1; if (ICED1EF5C0E5400F7869E1C674AE21DA6 > 1) IC52F3B77F7E45A74323561D6A6F6028A
<= 4'hf; end end I962095C6760357B792D0CD1278B21AF5 : begin I670A86ADD4DA92DA04F0354154D50812 <= 1'b1; if (IF4B2F356412545C21578876129150C2F )
I77B1E95A01761A9A5D153F6B403BCE8E <= {I2E664E814B6AA2CBCE57FBCE2A354435 , {14{1'b0}}, ICED1EF5C0E5400F7869E1C674AE21DA6 };
else I77B1E95A01761A9A5D153F6B403BCE8E <= {IEC10F95DD42CAF869EFB03BDF59BE8EB , {14{1'b0}}, ICED1EF5C0E5400F7869E1C674AE21DA6 };
end I9C2516A2CE92B199562345D5833785B3 : begin I670A86ADD4DA92DA04F0354154D50812 <= 1'b1; I77B1E95A01761A9A5D153F6B403BCE8E
<= {IF17B1273FDE2637DBFCD3D142F80E5D5 , I44E00CA48D123AE945CB7C612A95BFE6 , I5FC6334EB24FE23F5733F744B8E73624 ,
{8{1'b0}}, IC52F3B77F7E45A74323561D6A6F6028A , I11FD35FED78BCB8861FACB9A1E3A4C35 }; end I8A8F7A096F2E5012EDBEBDDEB9EEE34E
: begin I670A86ADD4DA92DA04F0354154D50812 <= 1'b1; if (IF4B2F356412545C21578876129150C2F ) I77B1E95A01761A9A5D153F6B403BCE8E
<= {{I1FC9733A3AF352A0F0C16A9487D3136E {1'b0}}, IE48F23B4AE45A1E423AC11ED564DE4D8 [I5D4944FED2815A3ECA7288050D4CB542
- 1:20]}; else begin I11FD35FED78BCB8861FACB9A1E3A4C35 <= {4{1'b1}}; IFFBEF8AE96EE878792DDB3FCC731CB4B <= &IABB783BAEC6EC4928216CD800CAC26FC ;
I1E515C54DF69EFC5334ACB78A7F46488 <= 1'b0; I77B1E95A01761A9A5D153F6B403BCE8E <= {IE48F23B4AE45A1E423AC11ED564DE4D8 [19:0],
I83C959FA1B0FD40F9B8261F8DA6D2791 , {2{1'b0}}}; I83C959FA1B0FD40F9B8261F8DA6D2791 <= IABB783BAEC6EC4928216CD800CAC26FC ;
if (IFFBEF8AE96EE878792DDB3FCC731CB4B ) begin IE48F23B4AE45A1E423AC11ED564DE4D8 <= IE48F23B4AE45A1E423AC11ED564DE4D8
+ 1; end end end IC6B19C3976DC11C4C29F6DFCC51BB3CF : begin I11FD35FED78BCB8861FACB9A1E3A4C35 <= {4{1'b1}}; IFFBEF8AE96EE878792DDB3FCC731CB4B
<= &IABB783BAEC6EC4928216CD800CAC26FC ; I1E515C54DF69EFC5334ACB78A7F46488 <= 1'b0; I670A86ADD4DA92DA04F0354154D50812
<= 1'b1; I77B1E95A01761A9A5D153F6B403BCE8E <= {IE48F23B4AE45A1E423AC11ED564DE4D8 [19:0], I83C959FA1B0FD40F9B8261F8DA6D2791 ,
{2{1'b0}}}; I83C959FA1B0FD40F9B8261F8DA6D2791 <= IABB783BAEC6EC4928216CD800CAC26FC ; if (IFFBEF8AE96EE878792DDB3FCC731CB4B )
begin IE48F23B4AE45A1E423AC11ED564DE4D8 <= IE48F23B4AE45A1E423AC11ED564DE4D8 + 1; end end I11ABAF7FCD68013E37F52A8A41493B59
: begin I0B6ECB7D58876821FA73D9499B8DE015 [9:0] <= ICED1EF5C0E5400F7869E1C674AE21DA6 ; I0B6ECB7D58876821FA73D9499B8DE015 [10]
<= ~(|ICED1EF5C0E5400F7869E1C674AE21DA6 ); I5A09FE74EFC8C7CD279F9D32F0E4BF2A <= (I0DE270F6B1F18A35E6835C0695437A55 )
? ~I21AD57B50E491E60E17CBE10D72C4241 : 1'b0; ICED1EF5C0E5400F7869E1C674AE21DA6 <= 0; end IEA810C9EE9AC978D2DFB6A0C31191743
: begin IF9EE6A022EB9CA07758C3F88273952CB <= 1'b0; I8D181359467F27637239CDAEE8A2F45A <= ~I8D181359467F27637239CDAEE8A2F45A
| (I8D181359467F27637239CDAEE8A2F45A & ~I24C403550AE065D7D1B7266142886226 ); end default : begin end endcase end
end endmodule 
  `timescale 1 ns / 1 ps
module I96EF4C28535915F06C7CA4A3F14655BA # (parameter I7292F55C07BFD7FB8A60D29FFC186275 = 32, parameter IDD54D6BED81F43FAE3E38E047FDC453C
= 4, parameter I61D0345D311EC6FFC08DDDECE5F6127A = 256 ) ( input wire ICCFB0F435B37370076102F325BC08D20 , input
wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire IC79EC9A9F373F4B71374BDF6EDD31DE6 , input wire I0B1584CC72F630A0464E5AEC9833BDC1 ,
input wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] I04BC24D2B6403E54A64DE9E6C9ABAA2B , input wire I22B24791BA0E7AA2C686B1B2D776C636 ,
output wire [$clog2(I61D0345D311EC6FFC08DDDECE5F6127A ) - 1:0] I89011D8BA1FC92A73CD875E098FE685C , output wire [I7292F55C07BFD7FB8A60D29FFC186275
- 1:0] I7D649F765882BD862315E777ABA5263F , output wire IEC0F7C6B7374DC46475F297465617F07 , output wire I705C64753A50CDA034B5ACB332D71768 ,
output wire [$clog2(I61D0345D311EC6FFC08DDDECE5F6127A + 1) - 1:0] I233E0C0C8E5150F0CD8258F276D93942 , output wire
IBE0D6810EBD63B5C428623C578CF6D3A , output wire I115E90220158F08B0465E99D7F2561D3 );  localparam I36A1B4EB5B5564A6ED7EA4D42856EFB4
= $clog2(I61D0345D311EC6FFC08DDDECE5F6127A ); localparam I2F8DC10449A1F24468235753BBC3B988 = $clog2(I61D0345D311EC6FFC08DDDECE5F6127A
+ 1); localparam IEF532EA44160288B0ED6812C670E4CDB = I7292F55C07BFD7FB8A60D29FFC186275 ; localparam IC123CC1DD854BDF232C22DA342143DED
= IDD54D6BED81F43FAE3E38E047FDC453C ; localparam I41D54753579217A07881641483914F62 = IDD54D6BED81F43FAE3E38E047FDC453C
+ 1;  reg [I36A1B4EB5B5564A6ED7EA4D42856EFB4 - 1:0] IF8FA22381AE98928C01C1A8EF2CB0DC6 ; reg [IEF532EA44160288B0ED6812C670E4CDB
- 1:0] I894F310391E6F0D90216157105D6D74E ; reg I4658BEBD88261965B56801558C4C44C4 ; reg I01F907CE74154BFFA0C1437099B21186 ;
reg [I2F8DC10449A1F24468235753BBC3B988 - 1:0] IE1A203A1BCBBA5F947F638C3DFB65BF8 ; reg ID079750A1760FEED5898B26A23289BAD ;
reg I28ACD74043EE392893ABFA4360DDCD11 ; wire I2FAC1854542B2B806297DF5B4733F9D2 ;  assign I89011D8BA1FC92A73CD875E098FE685C
= IF8FA22381AE98928C01C1A8EF2CB0DC6 ; assign I7D649F765882BD862315E777ABA5263F = I894F310391E6F0D90216157105D6D74E ;
assign IEC0F7C6B7374DC46475F297465617F07 = I4658BEBD88261965B56801558C4C44C4 ; assign I705C64753A50CDA034B5ACB332D71768
= I01F907CE74154BFFA0C1437099B21186 ; assign I233E0C0C8E5150F0CD8258F276D93942 = IE1A203A1BCBBA5F947F638C3DFB65BF8 ;
assign IBE0D6810EBD63B5C428623C578CF6D3A = ID079750A1760FEED5898B26A23289BAD ; assign I115E90220158F08B0465E99D7F2561D3
= I28ACD74043EE392893ABFA4360DDCD11 ;  assign I2FAC1854542B2B806297DF5B4733F9D2 = I22B24791BA0E7AA2C686B1B2D776C636
& ~ID079750A1760FEED5898B26A23289BAD ;  generate if (1'b1) begin : I50905559064282CED274D62360FCE175 reg [1:0] ICA80E74165E79AFA565A1A052BE49F09 ;
always @(posedge ICCFB0F435B37370076102F325BC08D20 or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin if (I9ED2A9117D3AEAF54CBA7AD69083BCB7
== 1'b0) begin IF8FA22381AE98928C01C1A8EF2CB0DC6 <= {I36A1B4EB5B5564A6ED7EA4D42856EFB4 {1'b0}}; I894F310391E6F0D90216157105D6D74E
<= {IEF532EA44160288B0ED6812C670E4CDB {1'b0}}; I4658BEBD88261965B56801558C4C44C4 <= 1'b0; I01F907CE74154BFFA0C1437099B21186
<= 1'b0; IE1A203A1BCBBA5F947F638C3DFB65BF8 <= I61D0345D311EC6FFC08DDDECE5F6127A ; ID079750A1760FEED5898B26A23289BAD
<= 1'b0; I28ACD74043EE392893ABFA4360DDCD11 <= 1'b0; end else begin if (IC79EC9A9F373F4B71374BDF6EDD31DE6 == 1'b1)
begin IF8FA22381AE98928C01C1A8EF2CB0DC6 <= {I36A1B4EB5B5564A6ED7EA4D42856EFB4 {1'b0}}; I4658BEBD88261965B56801558C4C44C4
<= 1'b0; I01F907CE74154BFFA0C1437099B21186 <= 1'b0; IE1A203A1BCBBA5F947F638C3DFB65BF8 <= I61D0345D311EC6FFC08DDDECE5F6127A ;
ID079750A1760FEED5898B26A23289BAD <= 1'b0; I28ACD74043EE392893ABFA4360DDCD11 <= 1'b0; end else begin I894F310391E6F0D90216157105D6D74E
<= I04BC24D2B6403E54A64DE9E6C9ABAA2B ; I4658BEBD88261965B56801558C4C44C4 <= I2FAC1854542B2B806297DF5B4733F9D2 ;
 ICA80E74165E79AFA565A1A052BE49F09 = {I0B1584CC72F630A0464E5AEC9833BDC1 , I2FAC1854542B2B806297DF5B4733F9D2 }; case
(ICA80E74165E79AFA565A1A052BE49F09 ) 2'b01: begin I01F907CE74154BFFA0C1437099B21186 <= (IE1A203A1BCBBA5F947F638C3DFB65BF8
== I41D54753579217A07881641483914F62 ) ? 1'b1 : I01F907CE74154BFFA0C1437099B21186 ; ID079750A1760FEED5898B26A23289BAD
<= ID079750A1760FEED5898B26A23289BAD | ((IE1A203A1BCBBA5F947F638C3DFB65BF8 == 1) ? 1'b1 : 1'b0); IE1A203A1BCBBA5F947F638C3DFB65BF8
<= IE1A203A1BCBBA5F947F638C3DFB65BF8 - 1; I28ACD74043EE392893ABFA4360DDCD11 <= (IE1A203A1BCBBA5F947F638C3DFB65BF8
== 2) ? 1'b1 : 1'b0; end 2'b10: begin I01F907CE74154BFFA0C1437099B21186 <= (IE1A203A1BCBBA5F947F638C3DFB65BF8 ==
IC123CC1DD854BDF232C22DA342143DED ) ? 1'b0 : I01F907CE74154BFFA0C1437099B21186 ; ID079750A1760FEED5898B26A23289BAD
<= 1'b0; IE1A203A1BCBBA5F947F638C3DFB65BF8 <= IE1A203A1BCBBA5F947F638C3DFB65BF8 + 1; I28ACD74043EE392893ABFA4360DDCD11
<= ID079750A1760FEED5898B26A23289BAD ; end endcase  if (I4658BEBD88261965B56801558C4C44C4 == 1'b1) IF8FA22381AE98928C01C1A8EF2CB0DC6
<= IF8FA22381AE98928C01C1A8EF2CB0DC6 + 1; end  end  end  end  endgenerate endmodule 
  `timescale 1 ns / 1 ps
module I1BD3AAA735BEFCAF06645830338869BC # (parameter I7292F55C07BFD7FB8A60D29FFC186275 = 32, parameter I7AEDD61970E812FD2535263A0E289FED
= 1, parameter ID93CAA7BF31348EA47B29E962BD456C7 = 4, parameter I61D0345D311EC6FFC08DDDECE5F6127A = 256 ) ( input
wire ICCFB0F435B37370076102F325BC08D20 , input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire [I7292F55C07BFD7FB8A60D29FFC186275
- 1 :0] I688B8620C444AB35D6A730AC46B175A1 , input wire IABAA7CE13DD3247C0A46E596E072DF77 , input wire IC79EC9A9F373F4B71374BDF6EDD31DE6 ,
input wire IFF897FEF3F69926A750D8217ADD6AE1C , output wire [$clog2(I61D0345D311EC6FFC08DDDECE5F6127A ) - 1:0] I7740E93179670969593F64CBA98864D9 ,
output wire I4101AA5DCE3023BCC2878E56C3794CB9 , output wire I11CEFC90537A67CD1FF01400245362F2 , output wire [$clog2((I61D0345D311EC6FFC08DDDECE5F6127A
* I7AEDD61970E812FD2535263A0E289FED ) + 1) - 1:0] ID7FCE45A65ADDB17F91F73A1B506BB5B , output wire [(I7292F55C07BFD7FB8A60D29FFC186275
/ I7AEDD61970E812FD2535263A0E289FED ) - 1:0] I125028C7446331521D0434C10E8B0007 , output wire I8BB939FF2AFDE7B2A1E480DCB61CE354 ,
output wire I41C63F948E534C7ED9F2471A44C922B2 , output wire I07E2A2E89C25B45C36871FC0931EC8EF );  localparam I36A1B4EB5B5564A6ED7EA4D42856EFB4
= $clog2(I61D0345D311EC6FFC08DDDECE5F6127A ); localparam I2F8DC10449A1F24468235753BBC3B988 = $clog2((I61D0345D311EC6FFC08DDDECE5F6127A
* I7AEDD61970E812FD2535263A0E289FED ) + 1); localparam I7759FD946E09EDD0DA617BA3BBAD1501 = I7292F55C07BFD7FB8A60D29FFC186275 ;
localparam ICA69BDD92A8EBD43E1DF50545F98A859 = I7292F55C07BFD7FB8A60D29FFC186275 / I7AEDD61970E812FD2535263A0E289FED ;
localparam I1AF585FFD3730CB75D8EA561C736B279 = ID93CAA7BF31348EA47B29E962BD456C7 ; localparam IB011AB9176BFCCD54AFA433401B9CC28
= ID93CAA7BF31348EA47B29E962BD456C7 + 1;  reg [I7AEDD61970E812FD2535263A0E289FED - 1:0] I10F60E589450CD09FF7A498641DE26F8 ;
reg I5C932555D8570D3003C70AC0892028C4 ; reg I38F39AED09C0507E780D3D35EA7FA06B ; reg [$clog2(I61D0345D311EC6FFC08DDDECE5F6127A )
- 1:0] I3283453B42BD77672B8ACE724ACDA314 ; reg I3B1A460AD69AD5EDF9D4E82F6E592EB8 ; reg I4FD65DDA0EDE2F39B09EF91789B31572 ;
reg [I2F8DC10449A1F24468235753BBC3B988 - 1:0] IDDFF27981262750D43304A01A2EBF659 ; reg [I7759FD946E09EDD0DA617BA3BBAD1501
- 1:0] I134B7C80786213E899F61495BA54C91C ; reg I00CE0BA4F77A2426865D797055E4C98A ; reg I35183CF475A58579BF332D0E77390724 ;
reg I8D7A3AECB8ADA4CFC13C707E28410478 ; reg IF084E43DB15C8EAD595BFBCBAB450494 ; reg I12B0B530CC957C3C059E79DA5211C283 ;
reg IFF286C818F68AC994E321B59884941FB ; wire [I7AEDD61970E812FD2535263A0E289FED - 1:0] IFF55929DAA63D5FAF40146769682E132 ;
wire I80D1B5313BBC5E22EAF77E255BDD847C ; wire IE699196B4C15D3DA4E93B2D4706C1C91 ; wire I09E9FB915D84D8A61BAF292FB1BDFA78 ;
 assign I7740E93179670969593F64CBA98864D9 = I3283453B42BD77672B8ACE724ACDA314 ; assign I4101AA5DCE3023BCC2878E56C3794CB9
= I38F39AED09C0507E780D3D35EA7FA06B ; assign I11CEFC90537A67CD1FF01400245362F2 = I4FD65DDA0EDE2F39B09EF91789B31572 ;
assign ID7FCE45A65ADDB17F91F73A1B506BB5B = IDDFF27981262750D43304A01A2EBF659 ; assign I125028C7446331521D0434C10E8B0007
= I134B7C80786213E899F61495BA54C91C [ICA69BDD92A8EBD43E1DF50545F98A859 - 1:0]; assign I8BB939FF2AFDE7B2A1E480DCB61CE354
= I00CE0BA4F77A2426865D797055E4C98A ; assign I41C63F948E534C7ED9F2471A44C922B2 = I35183CF475A58579BF332D0E77390724 ;
assign I07E2A2E89C25B45C36871FC0931EC8EF = IF084E43DB15C8EAD595BFBCBAB450494 ;  assign I80D1B5313BBC5E22EAF77E255BDD847C
= I10F60E589450CD09FF7A498641DE26F8 [0]; assign I09E9FB915D84D8A61BAF292FB1BDFA78 = IFF897FEF3F69926A750D8217ADD6AE1C
& ~I00CE0BA4F77A2426865D797055E4C98A & ~I8D7A3AECB8ADA4CFC13C707E28410478 ; generate if (I7AEDD61970E812FD2535263A0E289FED
== 1) begin assign IFF55929DAA63D5FAF40146769682E132 = 1'b1; assign IE699196B4C15D3DA4E93B2D4706C1C91 = I09E9FB915D84D8A61BAF292FB1BDFA78 ;
end else begin assign IFF55929DAA63D5FAF40146769682E132 = {I10F60E589450CD09FF7A498641DE26F8 [I7AEDD61970E812FD2535263A0E289FED
- 2:0], I10F60E589450CD09FF7A498641DE26F8 [I7AEDD61970E812FD2535263A0E289FED - 1]}; assign IE699196B4C15D3DA4E93B2D4706C1C91
= I09E9FB915D84D8A61BAF292FB1BDFA78 & I80D1B5313BBC5E22EAF77E255BDD847C ; end endgenerate  generate if (1'b1) begin :
I50905559064282CED274D62360FCE175 reg [1:0] I102EDFAABB65014FC78C55AF4345F765 ; always @(posedge ICCFB0F435B37370076102F325BC08D20
or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin if (I9ED2A9117D3AEAF54CBA7AD69083BCB7 == 1'b0) begin I10F60E589450CD09FF7A498641DE26F8
<= 1; I5C932555D8570D3003C70AC0892028C4 <= 1'b0; I38F39AED09C0507E780D3D35EA7FA06B <= 1'b0; I3283453B42BD77672B8ACE724ACDA314
<= {I36A1B4EB5B5564A6ED7EA4D42856EFB4 {1'b0}}; I3B1A460AD69AD5EDF9D4E82F6E592EB8 <= 1'b0; I4FD65DDA0EDE2F39B09EF91789B31572
<= 1'b0; IDDFF27981262750D43304A01A2EBF659 <= {I2F8DC10449A1F24468235753BBC3B988 {1'b0}}; I134B7C80786213E899F61495BA54C91C
<= {I7292F55C07BFD7FB8A60D29FFC186275 {1'b0}}; I00CE0BA4F77A2426865D797055E4C98A <= 1'b1; I35183CF475A58579BF332D0E77390724
<= 1'b0; I8D7A3AECB8ADA4CFC13C707E28410478 <= 1'b0; IF084E43DB15C8EAD595BFBCBAB450494 <= 1'b0; I12B0B530CC957C3C059E79DA5211C283
<= 1'b0; IFF286C818F68AC994E321B59884941FB <= 1'b0; end else begin if (IC79EC9A9F373F4B71374BDF6EDD31DE6 == 1'b1)
begin I10F60E589450CD09FF7A498641DE26F8 <= 1; I5C932555D8570D3003C70AC0892028C4 <= 1'b0; I38F39AED09C0507E780D3D35EA7FA06B
<= 1'b0; I3283453B42BD77672B8ACE724ACDA314 <= {I36A1B4EB5B5564A6ED7EA4D42856EFB4 {1'b0}}; I3B1A460AD69AD5EDF9D4E82F6E592EB8
<= 1'b0; I4FD65DDA0EDE2F39B09EF91789B31572 <= 1'b0; IDDFF27981262750D43304A01A2EBF659 <= {I2F8DC10449A1F24468235753BBC3B988 {1'b0}};
I00CE0BA4F77A2426865D797055E4C98A <= 1'b1; I35183CF475A58579BF332D0E77390724 <= 1'b0; I8D7A3AECB8ADA4CFC13C707E28410478
<= 1'b0; IF084E43DB15C8EAD595BFBCBAB450494 <= 1'b0; I12B0B530CC957C3C059E79DA5211C283 <= 1'b0; IFF286C818F68AC994E321B59884941FB
<= 1'b0; end else begin I5C932555D8570D3003C70AC0892028C4 <= I38F39AED09C0507E780D3D35EA7FA06B ; I38F39AED09C0507E780D3D35EA7FA06B
<= IE699196B4C15D3DA4E93B2D4706C1C91 ; I3B1A460AD69AD5EDF9D4E82F6E592EB8 <= IFF286C818F68AC994E321B59884941FB ;
I8D7A3AECB8ADA4CFC13C707E28410478 <= I09E9FB915D84D8A61BAF292FB1BDFA78 & I35183CF475A58579BF332D0E77390724 ; IF084E43DB15C8EAD595BFBCBAB450494
<= I12B0B530CC957C3C059E79DA5211C283 ; I12B0B530CC957C3C059E79DA5211C283 <= IFF286C818F68AC994E321B59884941FB ;
IFF286C818F68AC994E321B59884941FB <= I09E9FB915D84D8A61BAF292FB1BDFA78 ;  I102EDFAABB65014FC78C55AF4345F765 = {I09E9FB915D84D8A61BAF292FB1BDFA78 ,
IABAA7CE13DD3247C0A46E596E072DF77 }; case (I102EDFAABB65014FC78C55AF4345F765 ) 2'b01: begin I4FD65DDA0EDE2F39B09EF91789B31572
<= (IDDFF27981262750D43304A01A2EBF659 == I1AF585FFD3730CB75D8EA561C736B279 ) ? 1'b0 : I4FD65DDA0EDE2F39B09EF91789B31572 ;
I00CE0BA4F77A2426865D797055E4C98A <= 1'b0; IDDFF27981262750D43304A01A2EBF659 <= IDDFF27981262750D43304A01A2EBF659
+ I7AEDD61970E812FD2535263A0E289FED ; I35183CF475A58579BF332D0E77390724 <= (I7AEDD61970E812FD2535263A0E289FED ==
1) ? I00CE0BA4F77A2426865D797055E4C98A : 1'b0; end 2'b10: begin I4FD65DDA0EDE2F39B09EF91789B31572 <= (IDDFF27981262750D43304A01A2EBF659
== IB011AB9176BFCCD54AFA433401B9CC28 ) ? 1'b1 : I4FD65DDA0EDE2F39B09EF91789B31572 ; I00CE0BA4F77A2426865D797055E4C98A
<= I00CE0BA4F77A2426865D797055E4C98A | ((IDDFF27981262750D43304A01A2EBF659 == 1) ? 1'b1 : 1'b0); IDDFF27981262750D43304A01A2EBF659
<= IDDFF27981262750D43304A01A2EBF659 - 1; I35183CF475A58579BF332D0E77390724 <= (IDDFF27981262750D43304A01A2EBF659
== 2) ? 1'b1 : 1'b0; end 2'b11: begin I4FD65DDA0EDE2F39B09EF91789B31572 <= (IDDFF27981262750D43304A01A2EBF659 ==
I1AF585FFD3730CB75D8EA561C736B279 ) ? 1'b0 : I4FD65DDA0EDE2F39B09EF91789B31572 ; I00CE0BA4F77A2426865D797055E4C98A
<= 1'b0; IDDFF27981262750D43304A01A2EBF659 <= IDDFF27981262750D43304A01A2EBF659 + I7AEDD61970E812FD2535263A0E289FED
- 1; I35183CF475A58579BF332D0E77390724 <= (I7AEDD61970E812FD2535263A0E289FED == 1) ? ((IDDFF27981262750D43304A01A2EBF659
< 2) ? 1'b1 : 1'b0) : 1'b0; end default : begin I4FD65DDA0EDE2F39B09EF91789B31572 <= (IDDFF27981262750D43304A01A2EBF659
> I1AF585FFD3730CB75D8EA561C736B279 ) ? 1'b0 : I4FD65DDA0EDE2F39B09EF91789B31572 ; end endcase  if (I09E9FB915D84D8A61BAF292FB1BDFA78 )
I10F60E589450CD09FF7A498641DE26F8 <= IFF55929DAA63D5FAF40146769682E132 ; if (I5C932555D8570D3003C70AC0892028C4 )
I134B7C80786213E899F61495BA54C91C <= I688B8620C444AB35D6A730AC46B175A1 ; else if (I12B0B530CC957C3C059E79DA5211C283 )
I134B7C80786213E899F61495BA54C91C <= I134B7C80786213E899F61495BA54C91C >> (I7292F55C07BFD7FB8A60D29FFC186275 / I7AEDD61970E812FD2535263A0E289FED );
if (I38F39AED09C0507E780D3D35EA7FA06B ) I3283453B42BD77672B8ACE724ACDA314 <= I3283453B42BD77672B8ACE724ACDA314 +
1; end  end  end  end  endgenerate endmodule 
  `timescale 1 ns / 1 ps 
module I7C908B0C1EFA5CDE82E200D3BD5B8C53 # (parameter I18A8F7BCDF4CFE45E8382D66696B93B7 = 32, parameter IEC7FBEDC8625E773B8F1C7C89E5DA8F5
= 32, parameter IB71844FFA3AB85FEF45EAB4D35395752 = 512, parameter ID93CAA7BF31348EA47B29E962BD456C7 = 4, parameter
IDD54D6BED81F43FAE3E38E047FDC453C = 4, parameter I66C185998F46A7148163982E39BCD296 = "ecp3" ) ( input wire ICCFB0F435B37370076102F325BC08D20 ,
input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire IC79EC9A9F373F4B71374BDF6EDD31DE6 , input wire I48D61F5A0B5732A58912433B42CD9D0C ,
input wire [I18A8F7BCDF4CFE45E8382D66696B93B7 - 1:0] I04BC24D2B6403E54A64DE9E6C9ABAA2B , input wire IE315CDCA06C9620D5C0AB966E553F0C3 ,
output wire I11CEFC90537A67CD1FF01400245362F2 , output wire [$clog2((IB71844FFA3AB85FEF45EAB4D35395752 * (I18A8F7BCDF4CFE45E8382D66696B93B7 /IEC7FBEDC8625E773B8F1C7C89E5DA8F5 ))
+ 1) - 1:0] ID7FCE45A65ADDB17F91F73A1B506BB5B , output wire [IEC7FBEDC8625E773B8F1C7C89E5DA8F5 - 1:0] I125028C7446331521D0434C10E8B0007 ,
output wire I8BB939FF2AFDE7B2A1E480DCB61CE354 , output wire I41C63F948E534C7ED9F2471A44C922B2 , output wire I585F74DE05DD9C1C7070D6B4F6E181C2 ,
output wire I705C64753A50CDA034B5ACB332D71768 , output wire [$clog2(IB71844FFA3AB85FEF45EAB4D35395752 + 1) - 1:0]
I233E0C0C8E5150F0CD8258F276D93942 , output wire IBE0D6810EBD63B5C428623C578CF6D3A , output wire I115E90220158F08B0465E99D7F2561D3
);  localparam integer IE689EC19D4579850341747BD948B8E13 = I18A8F7BCDF4CFE45E8382D66696B93B7 / IEC7FBEDC8625E773B8F1C7C89E5DA8F5 ;
localparam integer I36A1B4EB5B5564A6ED7EA4D42856EFB4 = $clog2(IB71844FFA3AB85FEF45EAB4D35395752 ); localparam integer
I10B3AA6E839D478A1B149EA76A709877 = $clog2((IB71844FFA3AB85FEF45EAB4D35395752 * IE689EC19D4579850341747BD948B8E13 )
+ 1); localparam integer IE44C9D896DB0E0ECE64756576EED291E = $clog2(IB71844FFA3AB85FEF45EAB4D35395752 + 1); localparam
integer IF35F7B506981B2912E2486B227CB8871 = I18A8F7BCDF4CFE45E8382D66696B93B7 ;  wire [I36A1B4EB5B5564A6ED7EA4D42856EFB4
- 1:0] I75F7F62682CC33814DFF2B42BD851138 ; wire [IF35F7B506981B2912E2486B227CB8871 - 1:0] I8D9230DCE0724CC26C83BD6735F82BAB ;
wire I23CE9BB6FEF8024599BED6E7C9651049 ; wire I0E620501249C5CFBF447631D04D33715 ; wire [IE44C9D896DB0E0ECE64756576EED291E
- 1:0] I1E2790529716BDA31237F724D6F3C1DA ; wire I366EB0B781FD462E1BDC374519E76C20 ; wire IF63FD497AC79A293EAC51C0F982F9AD3 ;
wire [IF35F7B506981B2912E2486B227CB8871 - 1:0] I2CA1A324143051A0AFDEFB54659C657C ; wire [I36A1B4EB5B5564A6ED7EA4D42856EFB4
- 1:0] IB1475FB78BB097760DDF42DB8F04AFD0 ; wire IF8CBD565485880D1C0FCE2A4735DD796 ; wire IB52CCB2066E610613DDC71BD9DE3C046 ;
wire [I10B3AA6E839D478A1B149EA76A709877 - 1:0] I47BF20B234CB874608E4590CFA0DBE88 ; wire [IEC7FBEDC8625E773B8F1C7C89E5DA8F5
- 1:0] I967C0730B7C51D10FE97AFAB45FC31E4 ; wire IC7D9CDE692E08DD4B11A11E68738CB84 ; wire IA2B3584ECAB66E30B2B682D338F5CBA2 ;
wire I58AD4501D8BDFF58B28021F1FEDF600E ; wire I4AE98FF3DA4D5A5EE68F8A14D9D781F4 ;  assign I11CEFC90537A67CD1FF01400245362F2
= IB52CCB2066E610613DDC71BD9DE3C046 ; assign ID7FCE45A65ADDB17F91F73A1B506BB5B = I47BF20B234CB874608E4590CFA0DBE88 ;
assign I125028C7446331521D0434C10E8B0007 = I967C0730B7C51D10FE97AFAB45FC31E4 ; assign I8BB939FF2AFDE7B2A1E480DCB61CE354
= IC7D9CDE692E08DD4B11A11E68738CB84 ; assign I41C63F948E534C7ED9F2471A44C922B2 = IA2B3584ECAB66E30B2B682D338F5CBA2 ;
assign I585F74DE05DD9C1C7070D6B4F6E181C2 = I58AD4501D8BDFF58B28021F1FEDF600E ; assign I705C64753A50CDA034B5ACB332D71768
= I0E620501249C5CFBF447631D04D33715 ; assign I233E0C0C8E5150F0CD8258F276D93942 = I1E2790529716BDA31237F724D6F3C1DA ;
assign IBE0D6810EBD63B5C428623C578CF6D3A = I366EB0B781FD462E1BDC374519E76C20 ; assign I115E90220158F08B0465E99D7F2561D3
= IF63FD497AC79A293EAC51C0F982F9AD3 ;  assign I4AE98FF3DA4D5A5EE68F8A14D9D781F4 = ~I9ED2A9117D3AEAF54CBA7AD69083BCB7 ;
 I96EF4C28535915F06C7CA4A3F14655BA # ( .I7292F55C07BFD7FB8A60D29FFC186275 (I18A8F7BCDF4CFE45E8382D66696B93B7 ),
.IDD54D6BED81F43FAE3E38E047FDC453C (IDD54D6BED81F43FAE3E38E047FDC453C ), .I61D0345D311EC6FFC08DDDECE5F6127A (IB71844FFA3AB85FEF45EAB4D35395752 )
) I3133954E82C8A894470E1336CCBC8F15 ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .IC79EC9A9F373F4B71374BDF6EDD31DE6 (IC79EC9A9F373F4B71374BDF6EDD31DE6 ), .I0B1584CC72F630A0464E5AEC9833BDC1
(IF8CBD565485880D1C0FCE2A4735DD796 ), .I04BC24D2B6403E54A64DE9E6C9ABAA2B (I04BC24D2B6403E54A64DE9E6C9ABAA2B ), .I22B24791BA0E7AA2C686B1B2D776C636
(IE315CDCA06C9620D5C0AB966E553F0C3 ), .I89011D8BA1FC92A73CD875E098FE685C (I75F7F62682CC33814DFF2B42BD851138 ), .I7D649F765882BD862315E777ABA5263F
(I8D9230DCE0724CC26C83BD6735F82BAB ), .IEC0F7C6B7374DC46475F297465617F07 (I23CE9BB6FEF8024599BED6E7C9651049 ), .I705C64753A50CDA034B5ACB332D71768
(I0E620501249C5CFBF447631D04D33715 ), .I233E0C0C8E5150F0CD8258F276D93942 (I1E2790529716BDA31237F724D6F3C1DA ), .IBE0D6810EBD63B5C428623C578CF6D3A
(I366EB0B781FD462E1BDC374519E76C20 ), .I115E90220158F08B0465E99D7F2561D3 (IF63FD497AC79A293EAC51C0F982F9AD3 ) );
pmi_ram_dp # ( .pmi_wr_addr_depth (IB71844FFA3AB85FEF45EAB4D35395752 ), .pmi_wr_addr_width (I36A1B4EB5B5564A6ED7EA4D42856EFB4 ),
.pmi_wr_data_width (IF35F7B506981B2912E2486B227CB8871 ), .pmi_rd_addr_depth (IB71844FFA3AB85FEF45EAB4D35395752 ),
.pmi_rd_addr_width (I36A1B4EB5B5564A6ED7EA4D42856EFB4 ), .pmi_rd_data_width (IF35F7B506981B2912E2486B227CB8871 ),
.pmi_regmode ("reg"), .pmi_family (I66C185998F46A7148163982E39BCD296 ), .module_type ("pmi_ram_dp") ) I32900CECD80193336B4F376406D5DFF6
( .Data (I8D9230DCE0724CC26C83BD6735F82BAB ), .RdAddress (IB1475FB78BB097760DDF42DB8F04AFD0 ), .RdClockEn (1'b1),
.RdClock (ICCFB0F435B37370076102F325BC08D20 ), .Reset (I4AE98FF3DA4D5A5EE68F8A14D9D781F4 ), .WE (I23CE9BB6FEF8024599BED6E7C9651049 ),
.WrAddress (I75F7F62682CC33814DFF2B42BD851138 ), .WrClockEn (1'b1), .WrClock (ICCFB0F435B37370076102F325BC08D20 ),
.Q (I2CA1A324143051A0AFDEFB54659C657C ) ); I1BD3AAA735BEFCAF06645830338869BC # ( .I7292F55C07BFD7FB8A60D29FFC186275
(IF35F7B506981B2912E2486B227CB8871 ), .I7AEDD61970E812FD2535263A0E289FED (IE689EC19D4579850341747BD948B8E13 ), .ID93CAA7BF31348EA47B29E962BD456C7
(ID93CAA7BF31348EA47B29E962BD456C7 ), .I61D0345D311EC6FFC08DDDECE5F6127A (IB71844FFA3AB85FEF45EAB4D35395752 ) )
I306E1714C5A033192CADB7DE24CB682F ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .I688B8620C444AB35D6A730AC46B175A1 (I2CA1A324143051A0AFDEFB54659C657C ), .IABAA7CE13DD3247C0A46E596E072DF77
(I23CE9BB6FEF8024599BED6E7C9651049 ), .IC79EC9A9F373F4B71374BDF6EDD31DE6 (IC79EC9A9F373F4B71374BDF6EDD31DE6 ), .IFF897FEF3F69926A750D8217ADD6AE1C
(I48D61F5A0B5732A58912433B42CD9D0C ), .I7740E93179670969593F64CBA98864D9 (IB1475FB78BB097760DDF42DB8F04AFD0 ), .I4101AA5DCE3023BCC2878E56C3794CB9
(IF8CBD565485880D1C0FCE2A4735DD796 ), .I11CEFC90537A67CD1FF01400245362F2 (IB52CCB2066E610613DDC71BD9DE3C046 ), .ID7FCE45A65ADDB17F91F73A1B506BB5B
(I47BF20B234CB874608E4590CFA0DBE88 ), .I125028C7446331521D0434C10E8B0007 (I967C0730B7C51D10FE97AFAB45FC31E4 ), .I8BB939FF2AFDE7B2A1E480DCB61CE354
(IC7D9CDE692E08DD4B11A11E68738CB84 ), .I41C63F948E534C7ED9F2471A44C922B2 (IA2B3584ECAB66E30B2B682D338F5CBA2 ), .I07E2A2E89C25B45C36871FC0931EC8EF
(I58AD4501D8BDFF58B28021F1FEDF600E ) ); endmodule 
 module ID81B7D29F9F1B2882EE754B639B67517 # (parameter I7292F55C07BFD7FB8A60D29FFC186275 = 32, parameter IC3CEA40E2663BA267FBD739EE37AFBE9
= 512, parameter IAB32DAC10CBDBE04FD5EDBF7A576CAF9 = 512, parameter IB941270487D75F8FAA82F3DF028B6FC6 = 32, parameter
IFB129920FFBFCFD17ADB3180F882E8E1 = 48, parameter I66C185998F46A7148163982E39BCD296 = "ecp3" ) ( input wire ICCFB0F435B37370076102F325BC08D20 ,
input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire [7:0] IC680604FB338D55088F12313CDF2B03E , input wire [7:0]
IF17B1273FDE2637DBFCD3D142F80E5D5 , input wire [4:0] I44E00CA48D123AE945CB7C612A95BFE6 , input wire [2:0] I6D124B4E6D5F74B43E94949DE1CF46AA ,
input wire [2:0] I5C266315A3CF63C3FE988BB363C59AA1 , input wire I3EEFAC16E2400143CD0547F03531871C , input wire [IB941270487D75F8FAA82F3DF028B6FC6
- 1:0] I77DB6FE5680F7C0F4CCBA7F787115DDC , input wire I7AC0939DFAAFF38545186E63551C4452 , input wire [$clog2(IC3CEA40E2663BA267FBD739EE37AFBE9
+ 1) - 1:0] I10E4ABD5838C4A0B5C07B5A66417237D , input wire [$clog2(IAB32DAC10CBDBE04FD5EDBF7A576CAF9 + 1) - 1:0]
I3FF97406B3ED373B267711109A980AF9 , input wire I238A13C6F03704581F9A0A170F852FB4 , input wire I24C403550AE065D7D1B7266142886226 ,
input wire [IFB129920FFBFCFD17ADB3180F882E8E1 - 1:0] IDC6EA54AB52AEAD439CEF7521615AE1B , input wire [1:0] IC93EB5988EC451F72626A919FE396C61 ,
input wire [2:0] I6ED49B5BED4BA586759FFDCC7B3B7FF8 , input wire [7:0] I8E2F7CF6E50B95A483351A1836EB23AC , input
wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] I506D2FCB600E0189274870B654E65B64 , input wire [(I7292F55C07BFD7FB8A60D29FFC186275
/ 8) - 1:0] I1304D1B0EBC59FFD53EF6CD7A8537E4D , input wire I141300E29D7EF4A0D8B71CB7469A7B90 , input wire IC3CC91D317012C130AC9E2A126F71C64 ,
output wire [7:0] I7244B3A041E4EF91034ED304D36B4585 , output wire IC3E8DB22A270F4E2527F04E7E81EFA46 , output wire
IAEC671D12B80E2CC6E3D591A98E27230 , output wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] IA449B4CEADDC750F5446E3B900C14AA4 ,
output wire IFA413F55A4E38AA4A08DC60DCCB7553D , output wire I80F26623B387879BCA3F00C252D0129E , output wire [I7292F55C07BFD7FB8A60D29FFC186275
- 1:0] IFC7E490A5AF630CDD63895FB063ABE29 , output wire IEBE9989B3828CC1007CD10E6FBB2E76C , output wire I270ED686C2EF2C1C8B5B55EC4A5AAE84 ,
output wire IDA581E8478C8224118EF4E6B8EE8DDFE , output wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] I197028CF3B48BF15266050E66E13618E
);  localparam IE689EC19D4579850341747BD948B8E13 = IB941270487D75F8FAA82F3DF028B6FC6 / I7292F55C07BFD7FB8A60D29FFC186275 ;
localparam I6E124E2BABBAC497C974A94D29ED12FC = I7292F55C07BFD7FB8A60D29FFC186275 + 1;  wire [I7292F55C07BFD7FB8A60D29FFC186275 :0]
I42F9B19010F4C94942CB94E791F5B0A9 ; wire [7:0] I87F28D40CF2E19071DAC2CDAAC18501C ; wire [I7292F55C07BFD7FB8A60D29FFC186275
- 1:0] I0D700DE75DB58CB1498D11283A1D77A7 ; wire I7854B88F802C995C2468B7FAFE7E4680 ; wire IA7FB195B05854B5C9ADC134E6CEBE08D ;
wire I946A0D4483815E7E307A41EF5381B701 ; wire IE1B01EE52E8AB35666CA6D0FABD8DBB1 ; wire I5A6EEF2AFC2D0087CE28647E5950B7CD ;
wire I926EE9E5DB3F9321A6B286A451956E50 ; wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] I33241BB8F0FE626DE77345DEFE520975 ;
wire I8700EBE0E79B75823FD324C970684A6E ; wire IBB132FFAD30E399C86E32456EFA05229 ; wire [I7292F55C07BFD7FB8A60D29FFC186275
- 1:0] I395149947A0519460CDD6D133E28F6B9 ; wire IBABE4EF4D1FF12ED891304DB1676A43B ; wire I762EB11F447E9FE5C306D10B1D44F3D1 ;
wire I2FABB20E3D8A2178013BE94CDCF07251 ; wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] IDC4BF917DDF194B0E5BB9649E4071487 ;
wire [I7292F55C07BFD7FB8A60D29FFC186275 :0] I3332A83B1A159E66A80C07670C36A3BB ; wire IF04BEDCC6C3F0AE64FE5531D24835A27 ;
wire I47F5C1596C8EDF125D33B9CC7A68977B ; wire I4DDF7CB99428D62C1FB17E5C8FA42E6A ; wire I7DA036F5B0B44A1D5E3EB0237828A810 ;
wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] I0576740A3329B9B1A56E61643CACD3BB ; wire [$clog2(IAB32DAC10CBDBE04FD5EDBF7A576CAF9
+ 1) - 1:0] I7A3668BDA0446A1AEB107021676CD675 ;  assign I7244B3A041E4EF91034ED304D36B4585 = I87F28D40CF2E19071DAC2CDAAC18501C ;
assign IC3E8DB22A270F4E2527F04E7E81EFA46 = I5A6EEF2AFC2D0087CE28647E5950B7CD ; assign IAEC671D12B80E2CC6E3D591A98E27230
= I926EE9E5DB3F9321A6B286A451956E50 ; assign IA449B4CEADDC750F5446E3B900C14AA4 = I33241BB8F0FE626DE77345DEFE520975 ;
assign IFA413F55A4E38AA4A08DC60DCCB7553D = I8700EBE0E79B75823FD324C970684A6E ; assign I80F26623B387879BCA3F00C252D0129E
= IBB132FFAD30E399C86E32456EFA05229 ; assign IFC7E490A5AF630CDD63895FB063ABE29 = I395149947A0519460CDD6D133E28F6B9 ;
assign IEBE9989B3828CC1007CD10E6FBB2E76C = IBABE4EF4D1FF12ED891304DB1676A43B ; assign I270ED686C2EF2C1C8B5B55EC4A5AAE84
= I762EB11F447E9FE5C306D10B1D44F3D1 ; assign IDA581E8478C8224118EF4E6B8EE8DDFE = I2FABB20E3D8A2178013BE94CDCF07251 ;
assign I197028CF3B48BF15266050E66E13618E = IDC4BF917DDF194B0E5BB9649E4071487 ;  assign I42F9B19010F4C94942CB94E791F5B0A9
= {I7854B88F802C995C2468B7FAFE7E4680 , I0D700DE75DB58CB1498D11283A1D77A7 };  IC067A254D727EC6E4653DEA8E2C9ED79 #(
.I7292F55C07BFD7FB8A60D29FFC186275 (I7292F55C07BFD7FB8A60D29FFC186275 ), .I7AEDD61970E812FD2535263A0E289FED (IE689EC19D4579850341747BD948B8E13 ),
.I8B77F944A8EB2E113F742B8CB46E022C (IC3CEA40E2663BA267FBD739EE37AFBE9 ), .I5A1D0B7A4A119DC7A35D6729D171C67D (IAB32DAC10CBDBE04FD5EDBF7A576CAF9 ),
.ICFA9960F43620DB191960C5C79DBFAE6 (IAB32DAC10CBDBE04FD5EDBF7A576CAF9 ), .IFB129920FFBFCFD17ADB3180F882E8E1 (IFB129920FFBFCFD17ADB3180F882E8E1 )
) I2BFCA7961A4E4F9589575160D363B07A ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .IC680604FB338D55088F12313CDF2B03E (IC680604FB338D55088F12313CDF2B03E ), .IF17B1273FDE2637DBFCD3D142F80E5D5
(IF17B1273FDE2637DBFCD3D142F80E5D5 ), .I44E00CA48D123AE945CB7C612A95BFE6 (I44E00CA48D123AE945CB7C612A95BFE6 ), .I6D124B4E6D5F74B43E94949DE1CF46AA
(I6D124B4E6D5F74B43E94949DE1CF46AA ), .I5C266315A3CF63C3FE988BB363C59AA1 (I5C266315A3CF63C3FE988BB363C59AA1 ), .I8CE6978D396548B0C476A4C080ABF3CE
(I10E4ABD5838C4A0B5C07B5A66417237D ), .I879F5E0177BDD71945AEE80557DB31DC (I3332A83B1A159E66A80C07670C36A3BB [I7292F55C07BFD7FB8A60D29FFC186275
- 1:0]), .I3A0EE7E545E3C70F94B216D1405744A1 (I3332A83B1A159E66A80C07670C36A3BB [I7292F55C07BFD7FB8A60D29FFC186275 ]),
.I7B58D405D154321FAF23051CBA4F0967 (I7A3668BDA0446A1AEB107021676CD675 ), .I2FBCFC2E8A11BEE681E33A995F23A9F7 (IF04BEDCC6C3F0AE64FE5531D24835A27 ),
.I3EEFAC16E2400143CD0547F03531871C (I3EEFAC16E2400143CD0547F03531871C ), .I7AC0939DFAAFF38545186E63551C4452 (I7AC0939DFAAFF38545186E63551C4452 ),
.I9B878433B3D496FFA97B2BB22F930D6C (I47F5C1596C8EDF125D33B9CC7A68977B ), .I886DDC9EB90AFC1350E4197DB0F9F21D (I0576740A3329B9B1A56E61643CACD3BB ),
.IF63E3E7F031C0543230C8FA94864719C (I4DDF7CB99428D62C1FB17E5C8FA42E6A ), .I081430FC44E0C370F3B3B4FAFFC51A69 (I7DA036F5B0B44A1D5E3EB0237828A810 ),
.I3FF97406B3ED373B267711109A980AF9 (I3FF97406B3ED373B267711109A980AF9 ), .I238A13C6F03704581F9A0A170F852FB4 (I238A13C6F03704581F9A0A170F852FB4 ),
.I24C403550AE065D7D1B7266142886226 (I24C403550AE065D7D1B7266142886226 ), .IDC6EA54AB52AEAD439CEF7521615AE1B (IDC6EA54AB52AEAD439CEF7521615AE1B ),
.IC93EB5988EC451F72626A919FE396C61 (IC93EB5988EC451F72626A919FE396C61 ), .I6ED49B5BED4BA586759FFDCC7B3B7FF8 (I6ED49B5BED4BA586759FFDCC7B3B7FF8 ),
.I8E2F7CF6E50B95A483351A1836EB23AC (I8E2F7CF6E50B95A483351A1836EB23AC ), .I506D2FCB600E0189274870B654E65B64 (I506D2FCB600E0189274870B654E65B64 ),
.I1304D1B0EBC59FFD53EF6CD7A8537E4D (I1304D1B0EBC59FFD53EF6CD7A8537E4D ), .I141300E29D7EF4A0D8B71CB7469A7B90 (I141300E29D7EF4A0D8B71CB7469A7B90 ),
.IC3CC91D317012C130AC9E2A126F71C64 (IC3CC91D317012C130AC9E2A126F71C64 ), .I7244B3A041E4EF91034ED304D36B4585 (I87F28D40CF2E19071DAC2CDAAC18501C ),
.I37622C557C24CD88B10BAD5A6CB7A4F4 (I0D700DE75DB58CB1498D11283A1D77A7 ), .I1E2C39A87E460C8AD520B4134F92292F (I7854B88F802C995C2468B7FAFE7E4680 ),
.I406DAF97F28CB5044A320565BE60692E (IA7FB195B05854B5C9ADC134E6CEBE08D ), .ID24A83D781EA7F2CED8B0B12FADF20A5 (I946A0D4483815E7E307A41EF5381B701 ),
.IBADF395C0E67BC1FE7946C3D677241C4 (IE1B01EE52E8AB35666CA6D0FABD8DBB1 ), .IFB8B86C094497D5E859750490AB93CB4 ( ),
.IC3E8DB22A270F4E2527F04E7E81EFA46 (I5A6EEF2AFC2D0087CE28647E5950B7CD ), .IAEC671D12B80E2CC6E3D591A98E27230 (I926EE9E5DB3F9321A6B286A451956E50 ),
.IA449B4CEADDC750F5446E3B900C14AA4 (I33241BB8F0FE626DE77345DEFE520975 ), .IFA413F55A4E38AA4A08DC60DCCB7553D (I8700EBE0E79B75823FD324C970684A6E ),
.I80F26623B387879BCA3F00C252D0129E (IBB132FFAD30E399C86E32456EFA05229 ), .IFC7E490A5AF630CDD63895FB063ABE29 (I395149947A0519460CDD6D133E28F6B9 ),
.IEBE9989B3828CC1007CD10E6FBB2E76C (IBABE4EF4D1FF12ED891304DB1676A43B ), .I270ED686C2EF2C1C8B5B55EC4A5AAE84 (I762EB11F447E9FE5C306D10B1D44F3D1 ),
.IDA581E8478C8224118EF4E6B8EE8DDFE (I2FABB20E3D8A2178013BE94CDCF07251 ), .I197028CF3B48BF15266050E66E13618E (IDC4BF917DDF194B0E5BB9649E4071487 )
);  IF4FD65273243DC47A72869EEEA639DCD #( .I7292F55C07BFD7FB8A60D29FFC186275 (I6E124E2BABBAC497C974A94D29ED12FC ),
.IB71844FFA3AB85FEF45EAB4D35395752 (IAB32DAC10CBDBE04FD5EDBF7A576CAF9 ), .I66C185998F46A7148163982E39BCD296 (I66C185998F46A7148163982E39BCD296 )
) I7354CF0352544B8524D5654A5D14AD43 ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .IC79EC9A9F373F4B71374BDF6EDD31DE6 (1'b0), .I48D61F5A0B5732A58912433B42CD9D0C
(IA7FB195B05854B5C9ADC134E6CEBE08D ), .I04BC24D2B6403E54A64DE9E6C9ABAA2B (I42F9B19010F4C94942CB94E791F5B0A9 ), .IE315CDCA06C9620D5C0AB966E553F0C3
(I946A0D4483815E7E307A41EF5381B701 ), .I11CEFC90537A67CD1FF01400245362F2 (), .ID7FCE45A65ADDB17F91F73A1B506BB5B
(), .I125028C7446331521D0434C10E8B0007 (I3332A83B1A159E66A80C07670C36A3BB ), .I8BB939FF2AFDE7B2A1E480DCB61CE354
(), .I41C63F948E534C7ED9F2471A44C922B2 (), .I585F74DE05DD9C1C7070D6B4F6E181C2 (IF04BEDCC6C3F0AE64FE5531D24835A27 ),
.I705C64753A50CDA034B5ACB332D71768 (), .I233E0C0C8E5150F0CD8258F276D93942 (I7A3668BDA0446A1AEB107021676CD675 ),
.IBE0D6810EBD63B5C428623C578CF6D3A (), .I115E90220158F08B0465E99D7F2561D3 () );  I7C908B0C1EFA5CDE82E200D3BD5B8C53
#( .I18A8F7BCDF4CFE45E8382D66696B93B7 (IB941270487D75F8FAA82F3DF028B6FC6 ), .IEC7FBEDC8625E773B8F1C7C89E5DA8F5 (I7292F55C07BFD7FB8A60D29FFC186275 ),
.IB71844FFA3AB85FEF45EAB4D35395752 (IAB32DAC10CBDBE04FD5EDBF7A576CAF9 ), .I66C185998F46A7148163982E39BCD296 (I66C185998F46A7148163982E39BCD296 )
) IDD4356A81322E2CDA89609EEA437DC75 ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .IC79EC9A9F373F4B71374BDF6EDD31DE6 (1'b0), .I48D61F5A0B5732A58912433B42CD9D0C
(IE1B01EE52E8AB35666CA6D0FABD8DBB1 ), .I04BC24D2B6403E54A64DE9E6C9ABAA2B (I77DB6FE5680F7C0F4CCBA7F787115DDC ), .IE315CDCA06C9620D5C0AB966E553F0C3
(I7AC0939DFAAFF38545186E63551C4452 ), .I11CEFC90537A67CD1FF01400245362F2 (I47F5C1596C8EDF125D33B9CC7A68977B ), .ID7FCE45A65ADDB17F91F73A1B506BB5B
(), .I125028C7446331521D0434C10E8B0007 (I0576740A3329B9B1A56E61643CACD3BB ), .I8BB939FF2AFDE7B2A1E480DCB61CE354
(I4DDF7CB99428D62C1FB17E5C8FA42E6A ), .I41C63F948E534C7ED9F2471A44C922B2 (), .I585F74DE05DD9C1C7070D6B4F6E181C2
(I7DA036F5B0B44A1D5E3EB0237828A810 ), .I705C64753A50CDA034B5ACB332D71768 (), .I233E0C0C8E5150F0CD8258F276D93942
(), .IBE0D6810EBD63B5C428623C578CF6D3A (), .I115E90220158F08B0465E99D7F2561D3 () ); endmodule 
  module IF9CF184FC93B215506F993588C9E7793 #( parameter IA0A1D7DFDF0383A04E3B3C4C17E31A52 = "NONE", I1E00FE12AF273F059E9BCE9D0B8B6DCE
= 0, I41505CD673D5068189FBBD74B42776C5 = 0, I519B10D04CF8EB407876799C74F75633 = 1 ) ( input wire ICCFB0F435B37370076102F325BC08D20 ,
input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire [31:0] I9F8484FBCA62AC2BC8E1CB3333CC09DC , input wire
[31:0] I38F41A809C185C6FC2C37D7677D6013A , input wire I003A2455D9D9F27B56BE4B6A6E330845 , input wire I61583F0AD8ACE3D2B571B36EFC23311D ,
input wire I332C3203B01AAFA54A288D09DDEB7AFB , input wire I3D2849BFA4C1331FDDB8A39BF571CD91 , input wire [31:0]
I410A0939BF5AB6CE2A725DB6210E101F , input wire I22B24791BA0E7AA2C686B1B2D776C636 , output wire IAF378590D5A80382A321B73D17E05142 ,
output wire [31:0] IDCFC89CB36B3EFB6258338EC62FFDD79 ); `include "bar_reg_internals.v"
 reg I62799291AE8B63348A817ACCB8915B60 ; reg I8CD7C783B10692F81C0A4AE2406FA17C ; reg I356A069246FC6CDBCBD45DF848899082 ;
reg [31:0] I2A05666985F9532640F2423B1E7872D8 ; reg [31:0] I2D3AC641109F53FE7256D712A04790E2 ; reg I93FEA934E2F91A4D5E773376B9B26FED ;
reg I94914DEFD0BF8E6E975C4FECCB51F5B8 ; wire [5:0] I40F2C92F9483FEBACD49C34F556A2907 ; wire [3:0] IA1DF4C614A6FB93299EB3151A6E99586 ;
wire IC0D63F4CEDE2909E8A118A145BA3B6B9 ; wire [31:0] I5AD46C158BA68BFC32CD21A66C780D5E ; wire I87E5D05933CEDE6FA42E9E6B74C726DE ;
wire I1D7593F693FE0D78465004284368D454 ; wire [31:0] IBE741535D7456C7D7FC527AB8CFAD314 ;  assign IAF378590D5A80382A321B73D17E05142
= I1D7593F693FE0D78465004284368D454 ; assign IDCFC89CB36B3EFB6258338EC62FFDD79 = I2D3AC641109F53FE7256D712A04790E2
| {28'b0, IA1DF4C614A6FB93299EB3151A6E99586 };  generate begin if (I1E00FE12AF273F059E9BCE9D0B8B6DCE ) assign I87E5D05933CEDE6FA42E9E6B74C726DE
= 1'b1; else if (I41505CD673D5068189FBBD74B42776C5 ) begin if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "4") begin assign
I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 2; end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52
== "8") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 3; end
else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "16") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign
I40F2C92F9483FEBACD49C34F556A2907 = 4; end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "32") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE
= 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 5; end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "64") begin
assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 6; end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52
== "128") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 7; end
else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "256") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign
I40F2C92F9483FEBACD49C34F556A2907 = 8; end else begin assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b0; assign I40F2C92F9483FEBACD49C34F556A2907
= 0; end end else begin if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "128") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE
= 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 7; end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "256") begin
assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 8; end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52
== "512") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 9; end
else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "1K") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign
I40F2C92F9483FEBACD49C34F556A2907 = 10; end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "2K") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE
= 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 11; end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "4K") begin
assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 12; end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52
== "8K") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 13; end
else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "16K") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign
I40F2C92F9483FEBACD49C34F556A2907 = 14; end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "32K") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE
= 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 15; end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "64K")
begin assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 16; end else if
(IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "128K") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907
= 17; end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "256K") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE =
1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 18; end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "512K") begin
assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 19; end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52
== "1M") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 20; end
else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "2M") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign
I40F2C92F9483FEBACD49C34F556A2907 = 21; end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "4M") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE
= 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 22; end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "8M") begin
assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 23; end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52
== "16M") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 24;
end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "32M") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1;
assign I40F2C92F9483FEBACD49C34F556A2907 = 25; end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "64M") begin assign
I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 26; end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52
== "128M") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 27;
end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "256M") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1;
assign I40F2C92F9483FEBACD49C34F556A2907 = 28; end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "512M") begin assign
I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 29; end else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52
== "1G") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign I40F2C92F9483FEBACD49C34F556A2907 = 30; end
else if (IA0A1D7DFDF0383A04E3B3C4C17E31A52 == "2G") begin assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b1; assign
I40F2C92F9483FEBACD49C34F556A2907 = 31; end else begin assign I87E5D05933CEDE6FA42E9E6B74C726DE = 1'b0; assign I40F2C92F9483FEBACD49C34F556A2907
= 0; end end end endgenerate generate begin if (I1E00FE12AF273F059E9BCE9D0B8B6DCE ) assign IC0D63F4CEDE2909E8A118A145BA3B6B9
= 1'b1; else assign IC0D63F4CEDE2909E8A118A145BA3B6B9 = 1'b0; if (I1E00FE12AF273F059E9BCE9D0B8B6DCE ) assign IA1DF4C614A6FB93299EB3151A6E99586
= 4'b0; else assign IA1DF4C614A6FB93299EB3151A6E99586 = (I87E5D05933CEDE6FA42E9E6B74C726DE ) ? I6AD267363A4948AD568C784061BD44E6 (I41505CD673D5068189FBBD74B42776C5 ,
I1E00FE12AF273F059E9BCE9D0B8B6DCE , I519B10D04CF8EB407876799C74F75633 ) : 4'b0; assign I5AD46C158BA68BFC32CD21A66C780D5E
= I007A17D739E2006CB5D08DA8E8C1F04F (I40F2C92F9483FEBACD49C34F556A2907 , I41505CD673D5068189FBBD74B42776C5 , I1E00FE12AF273F059E9BCE9D0B8B6DCE );
end endgenerate  assign I1D7593F693FE0D78465004284368D454 = I356A069246FC6CDBCBD45DF848899082 & I93FEA934E2F91A4D5E773376B9B26FED
& I62799291AE8B63348A817ACCB8915B60 ; assign IBE741535D7456C7D7FC527AB8CFAD314 = I5AD46C158BA68BFC32CD21A66C780D5E
| {I2A05666985F9532640F2423B1E7872D8 [31:4], 4'b0};  always @(posedge ICCFB0F435B37370076102F325BC08D20 or negedge
I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin if (~I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin I62799291AE8B63348A817ACCB8915B60
<= 1'b0; I8CD7C783B10692F81C0A4AE2406FA17C <= 1'b0; I356A069246FC6CDBCBD45DF848899082 <= 1'b0; I2A05666985F9532640F2423B1E7872D8
<= 32'b0; I2D3AC641109F53FE7256D712A04790E2 <= 32'b0; I93FEA934E2F91A4D5E773376B9B26FED <= 1'b0; I94914DEFD0BF8E6E975C4FECCB51F5B8
<= 1'b0; end else begin I62799291AE8B63348A817ACCB8915B60 <= ((I9F8484FBCA62AC2BC8E1CB3333CC09DC & IBE741535D7456C7D7FC527AB8CFAD314 )
== (I2D3AC641109F53FE7256D712A04790E2 & IBE741535D7456C7D7FC527AB8CFAD314 )) ? 1'b1 : 1'b0; I356A069246FC6CDBCBD45DF848899082
<= I8CD7C783B10692F81C0A4AE2406FA17C & ((I003A2455D9D9F27B56BE4B6A6E330845 & IA1DF4C614A6FB93299EB3151A6E99586 [0])
| (I61583F0AD8ACE3D2B571B36EFC23311D & ~IA1DF4C614A6FB93299EB3151A6E99586 [0]) | (I61583F0AD8ACE3D2B571B36EFC23311D
& IC0D63F4CEDE2909E8A118A145BA3B6B9 )); I93FEA934E2F91A4D5E773376B9B26FED <= (I332C3203B01AAFA54A288D09DDEB7AFB
& IA1DF4C614A6FB93299EB3151A6E99586 [0]) | (I3D2849BFA4C1331FDDB8A39BF571CD91 & ~IA1DF4C614A6FB93299EB3151A6E99586 [0]
& ~IC0D63F4CEDE2909E8A118A145BA3B6B9 ) | (I3D2849BFA4C1331FDDB8A39BF571CD91 & IC0D63F4CEDE2909E8A118A145BA3B6B9 );
if (~I94914DEFD0BF8E6E975C4FECCB51F5B8 ) begin I2A05666985F9532640F2423B1E7872D8 <= I38F41A809C185C6FC2C37D7677D6013A ;
I94914DEFD0BF8E6E975C4FECCB51F5B8 <= 1'b1; end if (I22B24791BA0E7AA2C686B1B2D776C636 ) begin I8CD7C783B10692F81C0A4AE2406FA17C
<= I87E5D05933CEDE6FA42E9E6B74C726DE ; I2D3AC641109F53FE7256D712A04790E2 <= I410A0939BF5AB6CE2A725DB6210E101F &
IBE741535D7456C7D7FC527AB8CFAD314 ; end end end endmodule 
  module IDBAB269DB7AFDA96620B9B09A1C1D253 #( parameter I259BF2DBCEAAB39C062C08519379767E = 0, I2B0035459578DEB60AE2E24DF687E762
= 1, I2E554B9CAB59E598058B7921DA36D560 = "NONE", I86027F65FEA0494C8A49DAFE67EDAE13 = 0, ID3FF77989ABAC7B0FC1DE518FA7D21E6
= 1, IB04EEBB96EE0ED06EDBB60ACE60A4A93 = "NONE", ID022646F3454F5331B4174BB81BD0CF3 = 0 ) ( input wire ICCFB0F435B37370076102F325BC08D20 ,
input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire [31:0] I7195780B6CCA660A6833F98360035D81 , input wire
[31:0] I077B3A3A6F38E8073B18F35643BD4B02 , input wire [31:0] ICB680FEAB46B6D635CD9DD6BB49A6A20 , input wire [31:0]
I8FF768DAF4C56D1B2D217B2C02B6D4EC , input wire I003A2455D9D9F27B56BE4B6A6E330845 , input wire I61583F0AD8ACE3D2B571B36EFC23311D ,
input wire I332C3203B01AAFA54A288D09DDEB7AFB , input wire I3D2849BFA4C1331FDDB8A39BF571CD91 , input wire I94C1108CF14CB08354822C0EC9FFF090 ,
input wire I6E16E1B891ED18DC65EFF37952418F3C , input wire [31:0] I410A0939BF5AB6CE2A725DB6210E101F , input wire
I22B24791BA0E7AA2C686B1B2D776C636 , output wire [1:0] IAF378590D5A80382A321B73D17E05142 , output wire [31:0] IDCFC89CB36B3EFB6258338EC62FFDD79
);  wire IF95DF297621D7AF41FA0082F1A40C955 ; wire [31:0] I8CA75DECEF5DC240C5F341195D091889 ; wire IC5459C452507BEF54E88718AAB07CFA2 ;
wire [31:0] IC51CB268F59C6884F3B85925DA3F884B ; wire [31:0] I2610F1B6E08A8EF5DD0D052D30FCFA7B ; wire IA5052E8513A442F9E0B4D313BF0F3C24 ;
wire IDDCCC58C3FB71FE6E6701AA467ABE47B ; wire I65F18DE501DBD3CBB56BCEC8C26362EA ; wire I5E6DE37191562AC863CF1205F1C24780 ;
 assign IAF378590D5A80382A321B73D17E05142 = {IDDCCC58C3FB71FE6E6701AA467ABE47B , IA5052E8513A442F9E0B4D313BF0F3C24 };
assign IDCFC89CB36B3EFB6258338EC62FFDD79 = (I94C1108CF14CB08354822C0EC9FFF090 ) ? ((I6E16E1B891ED18DC65EFF37952418F3C )
? IC51CB268F59C6884F3B85925DA3F884B : I8CA75DECEF5DC240C5F341195D091889 ) : 32'b0;  assign I65F18DE501DBD3CBB56BCEC8C26362EA
= I22B24791BA0E7AA2C686B1B2D776C636 & I94C1108CF14CB08354822C0EC9FFF090 & I6E16E1B891ED18DC65EFF37952418F3C ; assign
I5E6DE37191562AC863CF1205F1C24780 = I22B24791BA0E7AA2C686B1B2D776C636 & I94C1108CF14CB08354822C0EC9FFF090 & ~I6E16E1B891ED18DC65EFF37952418F3C ;
 generate begin if (ID022646F3454F5331B4174BB81BD0CF3 ) begin assign I2610F1B6E08A8EF5DD0D052D30FCFA7B = I7195780B6CCA660A6833F98360035D81 ;
assign IA5052E8513A442F9E0B4D313BF0F3C24 = IF95DF297621D7AF41FA0082F1A40C955 & IC5459C452507BEF54E88718AAB07CFA2 ;
assign IDDCCC58C3FB71FE6E6701AA467ABE47B = 1'b0; end else begin assign I2610F1B6E08A8EF5DD0D052D30FCFA7B = I077B3A3A6F38E8073B18F35643BD4B02 ;
assign IA5052E8513A442F9E0B4D313BF0F3C24 = IF95DF297621D7AF41FA0082F1A40C955 ; assign IDDCCC58C3FB71FE6E6701AA467ABE47B
= IC5459C452507BEF54E88718AAB07CFA2 ; end end endgenerate  IF9CF184FC93B215506F993588C9E7793 #( .IA0A1D7DFDF0383A04E3B3C4C17E31A52
(I2E554B9CAB59E598058B7921DA36D560 ), .I1E00FE12AF273F059E9BCE9D0B8B6DCE (0), .I41505CD673D5068189FBBD74B42776C5
(I259BF2DBCEAAB39C062C08519379767E ), .I519B10D04CF8EB407876799C74F75633 (I2B0035459578DEB60AE2E24DF687E762 ) )
I33756A9C614D9965DC091F2B83660C43 ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .I9F8484FBCA62AC2BC8E1CB3333CC09DC (I077B3A3A6F38E8073B18F35643BD4B02 ), .I38F41A809C185C6FC2C37D7677D6013A
(ICB680FEAB46B6D635CD9DD6BB49A6A20 ), .I003A2455D9D9F27B56BE4B6A6E330845 (I003A2455D9D9F27B56BE4B6A6E330845 ), .I61583F0AD8ACE3D2B571B36EFC23311D
(I61583F0AD8ACE3D2B571B36EFC23311D ), .I332C3203B01AAFA54A288D09DDEB7AFB (I332C3203B01AAFA54A288D09DDEB7AFB ), .I3D2849BFA4C1331FDDB8A39BF571CD91
(I3D2849BFA4C1331FDDB8A39BF571CD91 ), .I410A0939BF5AB6CE2A725DB6210E101F (I410A0939BF5AB6CE2A725DB6210E101F ), .I22B24791BA0E7AA2C686B1B2D776C636
(I5E6DE37191562AC863CF1205F1C24780 ), .IAF378590D5A80382A321B73D17E05142 (IF95DF297621D7AF41FA0082F1A40C955 ), .IDCFC89CB36B3EFB6258338EC62FFDD79
(I8CA75DECEF5DC240C5F341195D091889 ) ); IF9CF184FC93B215506F993588C9E7793 #( .IA0A1D7DFDF0383A04E3B3C4C17E31A52
(IB04EEBB96EE0ED06EDBB60ACE60A4A93 ), .I1E00FE12AF273F059E9BCE9D0B8B6DCE (ID022646F3454F5331B4174BB81BD0CF3 ), .I41505CD673D5068189FBBD74B42776C5
(I86027F65FEA0494C8A49DAFE67EDAE13 ), .I519B10D04CF8EB407876799C74F75633 (ID3FF77989ABAC7B0FC1DE518FA7D21E6 ) )
IC2A14DD922AF115E3791DD3A0C8B3BE9 ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .I9F8484FBCA62AC2BC8E1CB3333CC09DC (I2610F1B6E08A8EF5DD0D052D30FCFA7B ), .I38F41A809C185C6FC2C37D7677D6013A
(I8FF768DAF4C56D1B2D217B2C02B6D4EC ), .I003A2455D9D9F27B56BE4B6A6E330845 (I003A2455D9D9F27B56BE4B6A6E330845 ), .I61583F0AD8ACE3D2B571B36EFC23311D
(I61583F0AD8ACE3D2B571B36EFC23311D ), .I332C3203B01AAFA54A288D09DDEB7AFB (I332C3203B01AAFA54A288D09DDEB7AFB ), .I3D2849BFA4C1331FDDB8A39BF571CD91
(I3D2849BFA4C1331FDDB8A39BF571CD91 ), .I410A0939BF5AB6CE2A725DB6210E101F (I410A0939BF5AB6CE2A725DB6210E101F ), .I22B24791BA0E7AA2C686B1B2D776C636
(I65F18DE501DBD3CBB56BCEC8C26362EA ), .IAF378590D5A80382A321B73D17E05142 (IC5459C452507BEF54E88718AAB07CFA2 ), .IDCFC89CB36B3EFB6258338EC62FFDD79
(IC51CB268F59C6884F3B85925DA3F884B ) ); endmodule 
  module I7649039BBE19689793FEE4FADDDEF1E8 #( parameter IFDFBBCC4A729BEC2BC4A96ABA6A686B0 = 0, I60C4892BECCA6E2B2FE143BD923A22CA
= 0, I614E1E615DEE042F64BC57A314245927 = 0, I2E554B9CAB59E598058B7921DA36D560 = "NONE", I259BF2DBCEAAB39C062C08519379767E
= 0, I2B0035459578DEB60AE2E24DF687E762 = 1, IB04EEBB96EE0ED06EDBB60ACE60A4A93 = "NONE", I86027F65FEA0494C8A49DAFE67EDAE13
= 0, ID3FF77989ABAC7B0FC1DE518FA7D21E6 = 1, IDD5BBB6DF3D487FCF2DA81CA8794849C = "NONE", I4E3CEE40D32239479A1163B2D85B5FA7
= 0, I41D8D6036479734032C1711509A67D83 = 1, I0AA7FFBF9C00DEF85FA40AFFAF675794 = "NONE", I6104B7636177E429318BE1C790C3CB49
= 0, I0D8F74FCCB77AD67CAB98890C8885156 = 1, IFB616CA07D005C26A9BA5823D543CCBD = "NONE", IA67F3F71E4F9434D68536978B81F91DA
= 0, IB6ECC5AF80982DE8999481CA0E9A481A = 1, I21FC0FBCD63A328488B305A90691197D = "NONE", I02E3D3076327F179BFEC2E663B0EAE70
= 0, I6D6B05AA28D91BF74A2607970B27F65D = 1 ) ( input wire ICCFB0F435B37370076102F325BC08D20 , input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 ,
input wire [31:0] I7195780B6CCA660A6833F98360035D81 , input wire [31:0] I077B3A3A6F38E8073B18F35643BD4B02 , input
wire I660A2BFC1099D715D966FB7D0E899778 , input wire I52BCA73A227659ABF278B7B041C2D33A , input wire I275F5F6495E251A9F1E0A46729B18393 ,
input wire [31:0] ICB680FEAB46B6D635CD9DD6BB49A6A20 , input wire [31:0] I8FF768DAF4C56D1B2D217B2C02B6D4EC , input
wire [31:0] I9E5E6E86745F53F982BC3862031A206B , input wire [31:0] I3AD72E1D6C16169DB8A27F1681293009 , input wire
[31:0] I0DE44F162EF92573C5DE1249527F6E9D , input wire [31:0] I2E9CC9AFC2E4742F852CB037CFC7E0A1 , input wire I003A2455D9D9F27B56BE4B6A6E330845 ,
input wire I61583F0AD8ACE3D2B571B36EFC23311D , input wire I332C3203B01AAFA54A288D09DDEB7AFB , input wire I3D2849BFA4C1331FDDB8A39BF571CD91 ,
input wire I6E16E1B891ED18DC65EFF37952418F3C , input wire [31:0] I410A0939BF5AB6CE2A725DB6210E101F , input wire
I22B24791BA0E7AA2C686B1B2D776C636 , output wire [5:0] IAF378590D5A80382A321B73D17E05142 , output wire [31:0] IDCFC89CB36B3EFB6258338EC62FFDD79
);  wire [1:0] IF95DF297621D7AF41FA0082F1A40C955 ; wire [31:0] I8CA75DECEF5DC240C5F341195D091889 ; wire [1:0] IC5459C452507BEF54E88718AAB07CFA2 ;
wire [31:0] IC51CB268F59C6884F3B85925DA3F884B ; wire [1:0] IDDF260B92ADEBC1228A3C40D8F02ABB2 ; wire [31:0] I8490321CB82DEFD9A157DA76A8FB74D1 ;
 assign IAF378590D5A80382A321B73D17E05142 = {IDDF260B92ADEBC1228A3C40D8F02ABB2 , IC5459C452507BEF54E88718AAB07CFA2 ,
IF95DF297621D7AF41FA0082F1A40C955 }; assign IDCFC89CB36B3EFB6258338EC62FFDD79 = I8CA75DECEF5DC240C5F341195D091889
| IC51CB268F59C6884F3B85925DA3F884B | I8490321CB82DEFD9A157DA76A8FB74D1 ;  IDBAB269DB7AFDA96620B9B09A1C1D253 #(
.I259BF2DBCEAAB39C062C08519379767E (I259BF2DBCEAAB39C062C08519379767E ), .I2B0035459578DEB60AE2E24DF687E762 (I2B0035459578DEB60AE2E24DF687E762 ),
.I2E554B9CAB59E598058B7921DA36D560 (I2E554B9CAB59E598058B7921DA36D560 ), .I86027F65FEA0494C8A49DAFE67EDAE13 (I86027F65FEA0494C8A49DAFE67EDAE13 ),
.ID3FF77989ABAC7B0FC1DE518FA7D21E6 (ID3FF77989ABAC7B0FC1DE518FA7D21E6 ), .IB04EEBB96EE0ED06EDBB60ACE60A4A93 (IB04EEBB96EE0ED06EDBB60ACE60A4A93 ),
.ID022646F3454F5331B4174BB81BD0CF3 (IFDFBBCC4A729BEC2BC4A96ABA6A686B0 ) ) I84BC79E638D11CEBD5CE37CCD54B92DA ( .ICCFB0F435B37370076102F325BC08D20
(ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .I7195780B6CCA660A6833F98360035D81
(I7195780B6CCA660A6833F98360035D81 ), .I077B3A3A6F38E8073B18F35643BD4B02 (I077B3A3A6F38E8073B18F35643BD4B02 ), .ICB680FEAB46B6D635CD9DD6BB49A6A20
(ICB680FEAB46B6D635CD9DD6BB49A6A20 ), .I8FF768DAF4C56D1B2D217B2C02B6D4EC (I8FF768DAF4C56D1B2D217B2C02B6D4EC ), .I003A2455D9D9F27B56BE4B6A6E330845
(I003A2455D9D9F27B56BE4B6A6E330845 ), .I61583F0AD8ACE3D2B571B36EFC23311D (I61583F0AD8ACE3D2B571B36EFC23311D ), .I332C3203B01AAFA54A288D09DDEB7AFB
(I332C3203B01AAFA54A288D09DDEB7AFB ), .I3D2849BFA4C1331FDDB8A39BF571CD91 (I3D2849BFA4C1331FDDB8A39BF571CD91 ), .I94C1108CF14CB08354822C0EC9FFF090
(I660A2BFC1099D715D966FB7D0E899778 ), .I6E16E1B891ED18DC65EFF37952418F3C (I6E16E1B891ED18DC65EFF37952418F3C ), .I410A0939BF5AB6CE2A725DB6210E101F
(I410A0939BF5AB6CE2A725DB6210E101F ), .I22B24791BA0E7AA2C686B1B2D776C636 (I22B24791BA0E7AA2C686B1B2D776C636 ), .IAF378590D5A80382A321B73D17E05142
(IF95DF297621D7AF41FA0082F1A40C955 ), .IDCFC89CB36B3EFB6258338EC62FFDD79 (I8CA75DECEF5DC240C5F341195D091889 ) );
IDBAB269DB7AFDA96620B9B09A1C1D253 #( .I259BF2DBCEAAB39C062C08519379767E (I4E3CEE40D32239479A1163B2D85B5FA7 ), .I2B0035459578DEB60AE2E24DF687E762
(I41D8D6036479734032C1711509A67D83 ), .I2E554B9CAB59E598058B7921DA36D560 (IDD5BBB6DF3D487FCF2DA81CA8794849C ), .I86027F65FEA0494C8A49DAFE67EDAE13
(I6104B7636177E429318BE1C790C3CB49 ), .ID3FF77989ABAC7B0FC1DE518FA7D21E6 (I0D8F74FCCB77AD67CAB98890C8885156 ), .IB04EEBB96EE0ED06EDBB60ACE60A4A93
(I0AA7FFBF9C00DEF85FA40AFFAF675794 ), .ID022646F3454F5331B4174BB81BD0CF3 (I60C4892BECCA6E2B2FE143BD923A22CA ) )
ID9BF48059D807303419933BF13879F87 ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .I7195780B6CCA660A6833F98360035D81 (I7195780B6CCA660A6833F98360035D81 ), .I077B3A3A6F38E8073B18F35643BD4B02
(I077B3A3A6F38E8073B18F35643BD4B02 ), .ICB680FEAB46B6D635CD9DD6BB49A6A20 (I9E5E6E86745F53F982BC3862031A206B ), .I8FF768DAF4C56D1B2D217B2C02B6D4EC
(I3AD72E1D6C16169DB8A27F1681293009 ), .I003A2455D9D9F27B56BE4B6A6E330845 (I003A2455D9D9F27B56BE4B6A6E330845 ), .I61583F0AD8ACE3D2B571B36EFC23311D
(I61583F0AD8ACE3D2B571B36EFC23311D ), .I332C3203B01AAFA54A288D09DDEB7AFB (I332C3203B01AAFA54A288D09DDEB7AFB ), .I3D2849BFA4C1331FDDB8A39BF571CD91
(I3D2849BFA4C1331FDDB8A39BF571CD91 ), .I94C1108CF14CB08354822C0EC9FFF090 (I52BCA73A227659ABF278B7B041C2D33A ), .I6E16E1B891ED18DC65EFF37952418F3C
(I6E16E1B891ED18DC65EFF37952418F3C ), .I410A0939BF5AB6CE2A725DB6210E101F (I410A0939BF5AB6CE2A725DB6210E101F ), .I22B24791BA0E7AA2C686B1B2D776C636
(I22B24791BA0E7AA2C686B1B2D776C636 ), .IAF378590D5A80382A321B73D17E05142 (IC5459C452507BEF54E88718AAB07CFA2 ), .IDCFC89CB36B3EFB6258338EC62FFDD79
(IC51CB268F59C6884F3B85925DA3F884B ) ); IDBAB269DB7AFDA96620B9B09A1C1D253 #( .I259BF2DBCEAAB39C062C08519379767E
(IA67F3F71E4F9434D68536978B81F91DA ), .I2B0035459578DEB60AE2E24DF687E762 (IB6ECC5AF80982DE8999481CA0E9A481A ), .I2E554B9CAB59E598058B7921DA36D560
(IFB616CA07D005C26A9BA5823D543CCBD ), .I86027F65FEA0494C8A49DAFE67EDAE13 (I02E3D3076327F179BFEC2E663B0EAE70 ), .ID3FF77989ABAC7B0FC1DE518FA7D21E6
(I6D6B05AA28D91BF74A2607970B27F65D ), .IB04EEBB96EE0ED06EDBB60ACE60A4A93 (I21FC0FBCD63A328488B305A90691197D ), .ID022646F3454F5331B4174BB81BD0CF3
(I614E1E615DEE042F64BC57A314245927 ) ) I8143B277EB85DE1485C118E148D5A9A4 ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ),
.I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .I7195780B6CCA660A6833F98360035D81 (I7195780B6CCA660A6833F98360035D81 ),
.I077B3A3A6F38E8073B18F35643BD4B02 (I077B3A3A6F38E8073B18F35643BD4B02 ), .ICB680FEAB46B6D635CD9DD6BB49A6A20 (I0DE44F162EF92573C5DE1249527F6E9D ),
.I8FF768DAF4C56D1B2D217B2C02B6D4EC (I2E9CC9AFC2E4742F852CB037CFC7E0A1 ), .I003A2455D9D9F27B56BE4B6A6E330845 (I003A2455D9D9F27B56BE4B6A6E330845 ),
.I61583F0AD8ACE3D2B571B36EFC23311D (I61583F0AD8ACE3D2B571B36EFC23311D ), .I332C3203B01AAFA54A288D09DDEB7AFB (I332C3203B01AAFA54A288D09DDEB7AFB ),
.I3D2849BFA4C1331FDDB8A39BF571CD91 (I3D2849BFA4C1331FDDB8A39BF571CD91 ), .I94C1108CF14CB08354822C0EC9FFF090 (I275F5F6495E251A9F1E0A46729B18393 ),
.I6E16E1B891ED18DC65EFF37952418F3C (I6E16E1B891ED18DC65EFF37952418F3C ), .I410A0939BF5AB6CE2A725DB6210E101F (I410A0939BF5AB6CE2A725DB6210E101F ),
.I22B24791BA0E7AA2C686B1B2D776C636 (I22B24791BA0E7AA2C686B1B2D776C636 ), .IAF378590D5A80382A321B73D17E05142 (IDDF260B92ADEBC1228A3C40D8F02ABB2 ),
.IDCFC89CB36B3EFB6258338EC62FFDD79 (I8490321CB82DEFD9A157DA76A8FB74D1 ) ); endmodule 
  module ID6D6E4DEEE2F225D2FE2E68AEDBFADC7 #( parameter I9449A4DEE4C71770D9A5095574AED415 = 0, parameter [23:0]
I4700AD5A2ED246219F585C312B2124C9 = 24'h000000, parameter [15:0] IB2FE05230F3A440BAF4BE98DCA56829F = 16'h0000, parameter
[5:0] I28B2C4B454208AC784C97EA8274B9503 = 0, parameter I7F482C6D7FFF305AD90ABABC0457155E = "INTA", parameter IBDE0431C8F903800F409661F4F56FD80
= 0, parameter [7:0] IE0E04F5EA496E6FD62B9A6B66E33F418 = 8'h00, parameter [15:0] I060C01BCB8E6DC3D4B74BEFA66D56545
= 16'h0000, parameter [15:0] ID34BC6EE8891CF37121D63EE0EAD6385 = 16'h0000, parameter [15:0] I9831646508922ACBA52B47759E0BAD32
= 16'h0000 ) ( input wire ICCFB0F435B37370076102F325BC08D20 , input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input
wire I1C0271AD5E8E9E9164909E468AD0B212 , input wire I9119CE851F731CBC5834D0370CCA6908 , input wire [11:0] I3D49ADB3C231E0C52B4EE7C42AB0DF8B ,
input wire [3:0] IE789C637CC57CC8ECB73F88C9790C5E4 , input wire [31:0] I3C3096B9DAB1C65EA381C7E05B767FB3 , input
wire I684F27663FD8A3EFB4B2BC8B42792CD0 , input wire I7378609E0B803011E82F6C6ABE861625 , output wire ICF9D8FD31DFC7D20DAF939C6D75F1518 ,
output wire IE4B6DD43E04940631EF58BA04EA58997 , output wire I3A095084CDFDFA56A0E67616A78D3B25 , output wire I81CD7F184DF8D58A1F2324E975A6816C ,
output wire I83C4A4200EB2B3F6766D338284ECAAAF , output wire IDA2B8A1BA5BD091F8C569BAA1CE5FED0 , output wire I9AFDACCEB4D156D714A2B8E72990FDA6 ,
output wire [31:0] IB808853736ABE6034DB8E375F1F00E89 ); `include "pcisig_constants.v"
 reg IBA8C2E9643A807EAD24886E1C89ED4E1 ; reg I0F63B15A4DE014E215E96C5F2D0B868F ; reg IFFAF919E74B9E78C820C15ECD6D17DDA ;
reg ICD9C74250F3A28D2BD3FCC4428D777F7 ; reg I9B8138DCE156F7C31EB5914EF01F183C ; reg [7:0] I98A5F7A73018ADA8369DAA8753CA8782 ;
reg [15:0] I260136A9A24C25C95FB2C4050C40596A ; reg [31:0] I72E47AC634CDDC2338CBBD5642F81090 ; reg [7:0] I9AA568501293D14DB94CBECC5A62ABD4 ;
reg I768376B2A960E56A7A0E19E757611EE3 ; reg [15:0] I58CBAA0FEF77AA53C1962EF903B6E7BB ; wire [7:0] IA6F6E55416AAFD05DDA78F9841BC80B4 ;
wire [7:0] IE2D0FB5EB0F870B2171CF15DBF995185 ; wire [7:0] I3319191F6960A33CEA37C0BE3D18B87E ; wire [7:0] I27F3E9958336B5B55EC5DD89EBD32846 ;
wire [7:0] I699007EC5E66211A0130F7D3AB75EE12 ; wire [7:0] I9310DFCF28F8C33DD2AFB8C0D2CEFACD ; wire I2CA2FB392686EFC907D0D5C7FFF051AD ;
wire [11:0] IDF2D2EFCFCAA060A180881D81395C002 ;  assign IDA2B8A1BA5BD091F8C569BAA1CE5FED0 = IFFAF919E74B9E78C820C15ECD6D17DDA ;
assign I9AFDACCEB4D156D714A2B8E72990FDA6 = ICD9C74250F3A28D2BD3FCC4428D777F7 ; assign ICF9D8FD31DFC7D20DAF939C6D75F1518
= IBA8C2E9643A807EAD24886E1C89ED4E1 ; assign IB808853736ABE6034DB8E375F1F00E89 = I7378609E0B803011E82F6C6ABE861625
? I72E47AC634CDDC2338CBBD5642F81090 : 32'b0;  generate if (I7F482C6D7FFF305AD90ABABC0457155E == "INTA") assign IE4B6DD43E04940631EF58BA04EA58997
= I768376B2A960E56A7A0E19E757611EE3 ; else assign IE4B6DD43E04940631EF58BA04EA58997 = 1'b0; if (I7F482C6D7FFF305AD90ABABC0457155E
== "INTB") assign I3A095084CDFDFA56A0E67616A78D3B25 = I768376B2A960E56A7A0E19E757611EE3 ; else assign I3A095084CDFDFA56A0E67616A78D3B25
= 1'b0; if (I7F482C6D7FFF305AD90ABABC0457155E == "INTC") assign I81CD7F184DF8D58A1F2324E975A6816C = I768376B2A960E56A7A0E19E757611EE3 ;
else assign I81CD7F184DF8D58A1F2324E975A6816C = 1'b0; if (I7F482C6D7FFF305AD90ABABC0457155E == "INTD") assign I83C4A4200EB2B3F6766D338284ECAAAF
= I768376B2A960E56A7A0E19E757611EE3 ; else assign I83C4A4200EB2B3F6766D338284ECAAAF = 1'b0; endgenerate  assign
I2CA2FB392686EFC907D0D5C7FFF051AD = I58CBAA0FEF77AA53C1962EF903B6E7BB [I07F7AABED30BAC0C4498CD527C624289 ] & ~I260136A9A24C25C95FB2C4050C40596A [I23FD9CC2F0EE3EAE050D08F50DC2BFA5 ]
& I9B8138DCE156F7C31EB5914EF01F183C & I0F63B15A4DE014E215E96C5F2D0B868F ; assign IDF2D2EFCFCAA060A180881D81395C002
= I3D49ADB3C231E0C52B4EE7C42AB0DF8B & 12'hffc;  generate begin assign IA6F6E55416AAFD05DDA78F9841BC80B4 = 8'h00;
assign IE2D0FB5EB0F870B2171CF15DBF995185 = I9449A4DEE4C71770D9A5095574AED415 ; if (I28B2C4B454208AC784C97EA8274B9503 )
if (I7F482C6D7FFF305AD90ABABC0457155E == "INTA") assign I27F3E9958336B5B55EC5DD89EBD32846 = I1A3B3F253A4CAA84340E1092DB0AD78B ;
else if (I7F482C6D7FFF305AD90ABABC0457155E == "INTB") assign I27F3E9958336B5B55EC5DD89EBD32846 = I496D2BA2FDE6A39BB367B7EC043A5D8A ;
else if (I7F482C6D7FFF305AD90ABABC0457155E == "INTC") assign I27F3E9958336B5B55EC5DD89EBD32846 = I0C9CD4F205090AE575352138FEB9E0B5 ;
else if (I7F482C6D7FFF305AD90ABABC0457155E == "INTD") assign I27F3E9958336B5B55EC5DD89EBD32846 = I5898D0798C075683D57F7DA612ED3F03 ;
else assign I27F3E9958336B5B55EC5DD89EBD32846 = 8'h00; else assign I27F3E9958336B5B55EC5DD89EBD32846 = 8'h00; if
(IBDE0431C8F903800F409661F4F56FD80 ) assign I3319191F6960A33CEA37C0BE3D18B87E = 8'h80; else assign I3319191F6960A33CEA37C0BE3D18B87E
= 8'h00; end endgenerate  always @(IDF2D2EFCFCAA060A180881D81395C002 or I7378609E0B803011E82F6C6ABE861625 ) begin
if (I7378609E0B803011E82F6C6ABE861625 ) case (IDF2D2EFCFCAA060A180881D81395C002 ) IF50924D3CD89C5522D937D4303186AAD
: I72E47AC634CDDC2338CBBD5642F81090 = {IB2FE05230F3A440BAF4BE98DCA56829F , I9831646508922ACBA52B47759E0BAD32 };
IE2B3CC108903457D70837BFC407A1BDB : I72E47AC634CDDC2338CBBD5642F81090 = {I58CBAA0FEF77AA53C1962EF903B6E7BB , I260136A9A24C25C95FB2C4050C40596A };
I6CDED12077023A013F4FB1192BA75334 : I72E47AC634CDDC2338CBBD5642F81090 = {I4700AD5A2ED246219F585C312B2124C9 , IE0E04F5EA496E6FD62B9A6B66E33F418 };
IF1FD22F074719F6000AB288899C22849 : I72E47AC634CDDC2338CBBD5642F81090 = {IA6F6E55416AAFD05DDA78F9841BC80B4 , I3319191F6960A33CEA37C0BE3D18B87E ,
8'h00, I98A5F7A73018ADA8369DAA8753CA8782 }; I14CB66CFC24FDF992E7D45E9D04A8A13 : I72E47AC634CDDC2338CBBD5642F81090
= {I060C01BCB8E6DC3D4B74BEFA66D56545 , ID34BC6EE8891CF37121D63EE0EAD6385 }; I6E0C77EC6D91F9E104E1B138A4446A8A :
I72E47AC634CDDC2338CBBD5642F81090 = { 24'h000000, IE2D0FB5EB0F870B2171CF15DBF995185 }; I9F4FDEC67E86458790E6BD886E959DE0
: I72E47AC634CDDC2338CBBD5642F81090 = { 16'h0000, I27F3E9958336B5B55EC5DD89EBD32846 , I9AA568501293D14DB94CBECC5A62ABD4 };
default : I72E47AC634CDDC2338CBBD5642F81090 = 32'b0; endcase else I72E47AC634CDDC2338CBBD5642F81090 = 32'b0; end
 always @(posedge ICCFB0F435B37370076102F325BC08D20 or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin if (~I9ED2A9117D3AEAF54CBA7AD69083BCB7 )
begin IBA8C2E9643A807EAD24886E1C89ED4E1 <= 1'b0; I0F63B15A4DE014E215E96C5F2D0B868F <= 1'b0; I768376B2A960E56A7A0E19E757611EE3
<= 1'b0; IFFAF919E74B9E78C820C15ECD6D17DDA <= 1'b0; ICD9C74250F3A28D2BD3FCC4428D777F7 <= 1'b0; I9B8138DCE156F7C31EB5914EF01F183C
<= 1'b0; I98A5F7A73018ADA8369DAA8753CA8782 <= 8'h00; I260136A9A24C25C95FB2C4050C40596A <= 16'h0000; I9AA568501293D14DB94CBECC5A62ABD4
<= 8'h00; I58CBAA0FEF77AA53C1962EF903B6E7BB <= 16'h0010; end else begin IBA8C2E9643A807EAD24886E1C89ED4E1 <= I260136A9A24C25C95FB2C4050C40596A [I146429BB43BA44B4E06CC733478550E1 ]
& I9B8138DCE156F7C31EB5914EF01F183C ; I0F63B15A4DE014E215E96C5F2D0B868F <= (|(I260136A9A24C25C95FB2C4050C40596A [1:0]))
? 1'b1 : 1'b0; I768376B2A960E56A7A0E19E757611EE3 <= I2CA2FB392686EFC907D0D5C7FFF051AD ; IFFAF919E74B9E78C820C15ECD6D17DDA
<= I260136A9A24C25C95FB2C4050C40596A [I9E02E8FD507F2B6814A8A105E77B80D5 ] & I9B8138DCE156F7C31EB5914EF01F183C ;
ICD9C74250F3A28D2BD3FCC4428D777F7 <= I260136A9A24C25C95FB2C4050C40596A [I245EA7B37D457CD05DEFB7F3E46EA478 ] & I9B8138DCE156F7C31EB5914EF01F183C ;
I9B8138DCE156F7C31EB5914EF01F183C <= I9119CE851F731CBC5834D0370CCA6908 ; I58CBAA0FEF77AA53C1962EF903B6E7BB [I07F7AABED30BAC0C4498CD527C624289 ]
<= I1C0271AD5E8E9E9164909E468AD0B212 ; if (I7378609E0B803011E82F6C6ABE861625 & I684F27663FD8A3EFB4B2BC8B42792CD0 )
case (IDF2D2EFCFCAA060A180881D81395C002 ) IE2B3CC108903457D70837BFC407A1BDB : begin if (IE789C637CC57CC8ECB73F88C9790C5E4 [0])
I260136A9A24C25C95FB2C4050C40596A [7:0] <= I3C3096B9DAB1C65EA381C7E05B767FB3 [7:0] & 8'h47; if (IE789C637CC57CC8ECB73F88C9790C5E4 [1])
I260136A9A24C25C95FB2C4050C40596A [15:8] <= I3C3096B9DAB1C65EA381C7E05B767FB3 [15:8] & 8'h05; end IF1FD22F074719F6000AB288899C22849
: begin if (IE789C637CC57CC8ECB73F88C9790C5E4 [0]) I98A5F7A73018ADA8369DAA8753CA8782 <= I3C3096B9DAB1C65EA381C7E05B767FB3 [7:0];
end I9F4FDEC67E86458790E6BD886E959DE0 : begin if (IE789C637CC57CC8ECB73F88C9790C5E4 [0]) I9AA568501293D14DB94CBECC5A62ABD4
<= I3C3096B9DAB1C65EA381C7E05B767FB3 [7:0]; end endcase end end endmodule 
  module IC3C2C92E294852CA4AE110FD59776962 #( parameter IF0D7F78B99E50997A728E3731A197225 = 0, I73ABD5619A9FB885445AC1E288EAF7F8
= 0 ) ( input wire ICCFB0F435B37370076102F325BC08D20 , input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire
IE145222FDBDC80109E12FA72D3D3C655 , input wire [2:0] I369BA2FFB5D41DF25F9BC3AB126D6607 , input wire I8E073ABA74C317770ABA5D59E6FA0BFF ,
input wire [31:0] I3C3096B9DAB1C65EA381C7E05B767FB3 , input wire [11:0] I438B8BD876741F9B46EB770E92F808B7 , input
wire I5FE75BE614D4F52DB327549B36203350 , input wire [31:0] I782B24592AE65A017A87162AE1B27668 , input wire [3:0]
I357B3043EDACE3EBECE8F54D79B9F90A , input wire I0AAD559CF33A5CBA597990658774FEB3 , input wire I923204A95D8CBB206587CF32BEDCF4EF ,
output wire I4A07557713C4283E634548A55A81AE55 , output wire IDF550B17734BF16B7E410B19BB31E276 , output wire [11:0]
I2E09014E801CDE025E646C14A7A88E8D , output wire [3:0] I095F5745EA5D8A16BF789BA5B07338AA , output wire [31:0] IB808853736ABE6034DB8E375F1F00E89 ,
output wire I14BCC8E29270920B2D04C15BCF409C2F , output wire I58DCF4F773FDA57377E940331963F6F2 , output wire I34D5C55E6A7E8D35B8981814BB90440B ,
output wire ID7CE65853F1A17B2A146805CE598364F , output wire I207147984DF21E60B2451E00D7A06100 , output wire I25F92BF03720992A727F6B9F19ACA644 ,
output wire I6A36AAB8630033974E1F982DFA8A6F7E , output wire I8B94BE4224AE909FF34FA01D95C810CE , output wire ID5CCD4858CB5CC1B2EDEC682C7DE5AAD ,
output wire [31:0] I6E43903839286F6F3DAB2A247E5C3D77 ); `include "pcisig_constants.v"
 reg I0DD988C25A5A5C0BBED3B2F0B83F6AE1 ; reg I30DDBB381375A42109F161AFFD0BA559 ; reg I05305DB38B053FE192F0B71598347D85 ;
reg I2D3F6195192E51E825219F43C080A709 ; reg [11:0] IC7779D4175ADF3F75C21392F9E824B6D ; reg ID564A30F71C7C1B827BA57264E89B21D ;
reg [31:0] I44109A75F9883AA09218902DA5B2CBB3 ; reg [31:0] I074FD9C5AE408613B3750B75A6125486 ; reg [3:0] I13C229A5BDE90D9F920D8F4D218106DE ;
reg I037773E6A298229B4A19627ABA272E81 ; reg I36FECBB048E15937DC767259CBABEDCB ; wire I895F10AA46CFA7CE62E6892D840FECE4 ;
wire I6533D1D0BB2CB6B5DD487B6DF8226F4B ; wire I6178D20A8C1F641D8C1EA99BA4484BA4 ; wire IE24FCD902B907F30C71F77BB6B81FBF7 ;
 assign I4A07557713C4283E634548A55A81AE55 = I0DD988C25A5A5C0BBED3B2F0B83F6AE1 ; assign IDF550B17734BF16B7E410B19BB31E276
= I30DDBB381375A42109F161AFFD0BA559 ; assign I2E09014E801CDE025E646C14A7A88E8D = (I6533D1D0BB2CB6B5DD487B6DF8226F4B )
? IC7779D4175ADF3F75C21392F9E824B6D : 12'b0; assign I095F5745EA5D8A16BF789BA5B07338AA = (IE24FCD902B907F30C71F77BB6B81FBF7 )
? I13C229A5BDE90D9F920D8F4D218106DE : 4'b0; assign IB808853736ABE6034DB8E375F1F00E89 = (IE24FCD902B907F30C71F77BB6B81FBF7 )
? I44109A75F9883AA09218902DA5B2CBB3 : 32'b0; assign I14BCC8E29270920B2D04C15BCF409C2F = (IE24FCD902B907F30C71F77BB6B81FBF7 )
? I36FECBB048E15937DC767259CBABEDCB : 1'b0; assign I58DCF4F773FDA57377E940331963F6F2 = ((IC7779D4175ADF3F75C21392F9E824B6D
== I59630A699E2E8DE4A02E477B2CE20A7D ) || (IC7779D4175ADF3F75C21392F9E824B6D == I4C0348AD8EE23C00D0A9F4C040509DD3 ))
? I6533D1D0BB2CB6B5DD487B6DF8226F4B : 1'b0; assign I34D5C55E6A7E8D35B8981814BB90440B = ((IC7779D4175ADF3F75C21392F9E824B6D
== I57D1D6FAFB22D1FFE8478966E395EF69 ) || (IC7779D4175ADF3F75C21392F9E824B6D == I132B6BD74FA99D570BBF433782EA41BE ))
? I6533D1D0BB2CB6B5DD487B6DF8226F4B : 1'b0; assign ID7CE65853F1A17B2A146805CE598364F = ((IC7779D4175ADF3F75C21392F9E824B6D
== IBB50DFD4A7725440E2A7F9205780698F ) || (IC7779D4175ADF3F75C21392F9E824B6D == I91282DABBD48120D1700BB2A213A5A33 ))
? I6533D1D0BB2CB6B5DD487B6DF8226F4B : 1'b0; assign I6A36AAB8630033974E1F982DFA8A6F7E = ((IC7779D4175ADF3F75C21392F9E824B6D
== I8125345218ED2F68A2205656CAD621A2 ) || (IC7779D4175ADF3F75C21392F9E824B6D == I9F1C08850EAFD27114AE21872A780597 ))
? I6533D1D0BB2CB6B5DD487B6DF8226F4B : 1'b0; assign I207147984DF21E60B2451E00D7A06100 = I895F10AA46CFA7CE62E6892D840FECE4 ;
assign I25F92BF03720992A727F6B9F19ACA644 = ((IC7779D4175ADF3F75C21392F9E824B6D >= IC8E275CE62D6604F5CC30E6E067A1EA0 )
&& (IC7779D4175ADF3F75C21392F9E824B6D < (IC8E275CE62D6604F5CC30E6E067A1EA0 + I5B58B630DCD4895F11E6244BDE0B377D )))
? I6533D1D0BB2CB6B5DD487B6DF8226F4B : 1'b0; assign I8B94BE4224AE909FF34FA01D95C810CE = ((IC7779D4175ADF3F75C21392F9E824B6D
< I59630A699E2E8DE4A02E477B2CE20A7D ) || ((IC7779D4175ADF3F75C21392F9E824B6D > I91282DABBD48120D1700BB2A213A5A33 )
&& (IC7779D4175ADF3F75C21392F9E824B6D < 12'h040))) ? I6533D1D0BB2CB6B5DD487B6DF8226F4B : 1'b0; assign ID5CCD4858CB5CC1B2EDEC682C7DE5AAD
= I2D3F6195192E51E825219F43C080A709 ; assign I6E43903839286F6F3DAB2A247E5C3D77 = I074FD9C5AE408613B3750B75A6125486 ;
 assign I6533D1D0BB2CB6B5DD487B6DF8226F4B = ID564A30F71C7C1B827BA57264E89B21D & I037773E6A298229B4A19627ABA272E81 ;
assign I6178D20A8C1F641D8C1EA99BA4484BA4 = ID564A30F71C7C1B827BA57264E89B21D & I037773E6A298229B4A19627ABA272E81
& ~I2D3F6195192E51E825219F43C080A709 ; assign IE24FCD902B907F30C71F77BB6B81FBF7 = I5FE75BE614D4F52DB327549B36203350
& I0AAD559CF33A5CBA597990658774FEB3 & I2D3F6195192E51E825219F43C080A709 ; generate if (IF0D7F78B99E50997A728E3731A197225 )
assign I895F10AA46CFA7CE62E6892D840FECE4 = ((IC7779D4175ADF3F75C21392F9E824B6D >= I43C945338ADA718C47F9AC36AE9ADB8A )
&& (IC7779D4175ADF3F75C21392F9E824B6D < (I43C945338ADA718C47F9AC36AE9ADB8A + I3BD1B3B7A6666C5993CC8BE2E2E17B9C )))
? I6533D1D0BB2CB6B5DD487B6DF8226F4B : 1'b0; else assign I895F10AA46CFA7CE62E6892D840FECE4 = 1'b0; endgenerate  always
@(posedge ICCFB0F435B37370076102F325BC08D20 or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin if (~I9ED2A9117D3AEAF54CBA7AD69083BCB7 )
begin I0DD988C25A5A5C0BBED3B2F0B83F6AE1 <= 1'b0; I30DDBB381375A42109F161AFFD0BA559 <= 1'b0; I05305DB38B053FE192F0B71598347D85
<= 1'b0; I2D3F6195192E51E825219F43C080A709 <= 1'b0; I074FD9C5AE408613B3750B75A6125486 <= 32'b0; IC7779D4175ADF3F75C21392F9E824B6D
<= 12'b0; ID564A30F71C7C1B827BA57264E89B21D <= 1'b0; I44109A75F9883AA09218902DA5B2CBB3 <= 32'b0; I13C229A5BDE90D9F920D8F4D218106DE
<= 4'b0; I037773E6A298229B4A19627ABA272E81 <= 1'b0; I36FECBB048E15937DC767259CBABEDCB <= 1'b0; end else begin I0DD988C25A5A5C0BBED3B2F0B83F6AE1
<= (I369BA2FFB5D41DF25F9BC3AB126D6607 == I73ABD5619A9FB885445AC1E288EAF7F8 ) ? IE145222FDBDC80109E12FA72D3D3C655
: 1'b0; I30DDBB381375A42109F161AFFD0BA559 <= I8E073ABA74C317770ABA5D59E6FA0BFF ; I05305DB38B053FE192F0B71598347D85
<= ID564A30F71C7C1B827BA57264E89B21D & I037773E6A298229B4A19627ABA272E81 & ~I36FECBB048E15937DC767259CBABEDCB &
~I2D3F6195192E51E825219F43C080A709 ; I2D3F6195192E51E825219F43C080A709 <= ((I5FE75BE614D4F52DB327549B36203350 &
I0AAD559CF33A5CBA597990658774FEB3 & I923204A95D8CBB206587CF32BEDCF4EF & ~I2D3F6195192E51E825219F43C080A709 ) | (ID564A30F71C7C1B827BA57264E89B21D
& I037773E6A298229B4A19627ABA272E81 & ~I36FECBB048E15937DC767259CBABEDCB & I6178D20A8C1F641D8C1EA99BA4484BA4 ))
& I0DD988C25A5A5C0BBED3B2F0B83F6AE1 ; I074FD9C5AE408613B3750B75A6125486 <= (I6178D20A8C1F641D8C1EA99BA4484BA4 )
? I3C3096B9DAB1C65EA381C7E05B767FB3 : 32'b0; IC7779D4175ADF3F75C21392F9E824B6D <= {I438B8BD876741F9B46EB770E92F808B7 [11:2],
2'b0}; ID564A30F71C7C1B827BA57264E89B21D <= I5FE75BE614D4F52DB327549B36203350 & ~I2D3F6195192E51E825219F43C080A709 ;
I44109A75F9883AA09218902DA5B2CBB3 <= I782B24592AE65A017A87162AE1B27668 ; I13C229A5BDE90D9F920D8F4D218106DE <= I357B3043EDACE3EBECE8F54D79B9F90A ;
I037773E6A298229B4A19627ABA272E81 <= I0AAD559CF33A5CBA597990658774FEB3 & ~I2D3F6195192E51E825219F43C080A709 ; I36FECBB048E15937DC767259CBABEDCB
<= I923204A95D8CBB206587CF32BEDCF4EF & ~I2D3F6195192E51E825219F43C080A709 ; end end endmodule 
 module ICD3F460CCA1DA6A6D1EAF48665780088 #( parameter I73ABD5619A9FB885445AC1E288EAF7F8 = 0 ) ( input wire ICCFB0F435B37370076102F325BC08D20 ,
input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire [7:0] I3C7A9FA839F554D8898020C4831479E2 , input wire [4:0]
I74A0936EE8FD1443A2C6745A4F3F6B5E , input wire [7:0] I691085C332A55972BA4126AE83875679 , input wire I1C0271AD5E8E9E9164909E468AD0B212 ,
input wire I56148DDDF284443347FFCF4F9C3BE61A , input wire I24C403550AE065D7D1B7266142886226 , output wire [31:0]
IFE4A8CBA73734C6F0F0A078027E053D4 , output wire ID7A2A8B1E9D92B60194D5FAFAAB15208 , output wire IF274FAF97F5BACD693913BB418717A9D ,
output wire ID95C13E7EE1CFE6A8743FF9E62C25873 , output wire [10:0] IC58E411F24D810EF60A7B8638ABCC0BB , output wire
I89CFFA73C7546481B72B0FB06D799AEE , output wire I270ED686C2EF2C1C8B5B55EC4A5AAE84 ); `include "pcisig_constants.v"
 localparam IBE3FC19439FEC0073D66B4DAC2FECC32 = 4'b0000, I310264643E51C96BF8FECF37C2EB7553 = 4'b0001, IA7E2C061B23F9C2D79751962637FF9F8
= 4'b0010, I0FBF38AB1DE3B938794F64EFEB6EEF04 = 4'b0011, I2512657214BD8CD9D7C9E46341FB6960 = 4'b0100, IA4F9276F2E3EF93B14F2B0FF3B2DDE74
= 4'b0101, I3AEAA310DC2EB1E6D2E2AB4DD0417BA2 = 4'b0110, I9CFCF3FC76F8BCD4AA7E722E67E01A89 = 4'b0111, IDA65D1282C0B7B2A86436F0450F882A3
= 4'b1000;  reg I37A362329A50BFF771D5547766A00B10 ; reg I2CA2FB392686EFC907D0D5C7FFF051AD ; reg IBE5A77ED6624B1E16464A1925007FB7C ;
reg [31:0] ID0A5ECECBEC8CE692F380DDF069E842F ; reg I1877CB8174894BB7A9732E91A1794AAA ; reg [3:0] I7E04E8229BE60B48AAE3E1EB6511163A ;
reg [3:0] ID22BB0550BCC1515614C8142FADDA171 ; reg I612E93B17FEB6E7AE6FD9448B52CA816 ; reg [10:0] I95FD0A1F8137860FD05FEA74508A613F ;
reg I09934DCB789133B6EE69ED6ABA942F05 ; reg I8D181359467F27637239CDAEE8A2F45A ; wire [2:0] IEAB12A55F034325A3F47B7F5B88B077D ;
wire I5EA9375131D29CCE63A1B4FB334D5BBD ;  assign IFE4A8CBA73734C6F0F0A078027E053D4 = ID0A5ECECBEC8CE692F380DDF069E842F ;
assign ID7A2A8B1E9D92B60194D5FAFAAB15208 = I1877CB8174894BB7A9732E91A1794AAA ; assign IF274FAF97F5BACD693913BB418717A9D
= I612E93B17FEB6E7AE6FD9448B52CA816 ; assign ID95C13E7EE1CFE6A8743FF9E62C25873 = (I7E04E8229BE60B48AAE3E1EB6511163A
== I310264643E51C96BF8FECF37C2EB7553 ) ? 1'b1 : 1'b0; assign IC58E411F24D810EF60A7B8638ABCC0BB = I95FD0A1F8137860FD05FEA74508A613F ;
assign I89CFFA73C7546481B72B0FB06D799AEE = I09934DCB789133B6EE69ED6ABA942F05 ; assign I270ED686C2EF2C1C8B5B55EC4A5AAE84
= I8D181359467F27637239CDAEE8A2F45A ;  assign I5EA9375131D29CCE63A1B4FB334D5BBD = (I7E04E8229BE60B48AAE3E1EB6511163A
== I9CFCF3FC76F8BCD4AA7E722E67E01A89 ) ? 1'b1 : 1'b0;  generate assign IEAB12A55F034325A3F47B7F5B88B077D = I73ABD5619A9FB885445AC1E288EAF7F8 ;
endgenerate  always @(I37A362329A50BFF771D5547766A00B10 or I7E04E8229BE60B48AAE3E1EB6511163A or I56148DDDF284443347FFCF4F9C3BE61A
or I24C403550AE065D7D1B7266142886226 ) begin ID22BB0550BCC1515614C8142FADDA171 = I7E04E8229BE60B48AAE3E1EB6511163A ;
case (I7E04E8229BE60B48AAE3E1EB6511163A ) IBE3FC19439FEC0073D66B4DAC2FECC32 : begin if (I37A362329A50BFF771D5547766A00B10 )
ID22BB0550BCC1515614C8142FADDA171 = I310264643E51C96BF8FECF37C2EB7553 ; end I310264643E51C96BF8FECF37C2EB7553 :
begin if (I56148DDDF284443347FFCF4F9C3BE61A ) ID22BB0550BCC1515614C8142FADDA171 = IA7E2C061B23F9C2D79751962637FF9F8 ;
end IA7E2C061B23F9C2D79751962637FF9F8 : begin ID22BB0550BCC1515614C8142FADDA171 = I0FBF38AB1DE3B938794F64EFEB6EEF04 ;
end I0FBF38AB1DE3B938794F64EFEB6EEF04 : begin ID22BB0550BCC1515614C8142FADDA171 = I2512657214BD8CD9D7C9E46341FB6960 ;
end I2512657214BD8CD9D7C9E46341FB6960 : begin ID22BB0550BCC1515614C8142FADDA171 = IA4F9276F2E3EF93B14F2B0FF3B2DDE74 ;
end IA4F9276F2E3EF93B14F2B0FF3B2DDE74 : begin ID22BB0550BCC1515614C8142FADDA171 = I3AEAA310DC2EB1E6D2E2AB4DD0417BA2 ;
end I3AEAA310DC2EB1E6D2E2AB4DD0417BA2 : begin ID22BB0550BCC1515614C8142FADDA171 = I9CFCF3FC76F8BCD4AA7E722E67E01A89 ;
end I9CFCF3FC76F8BCD4AA7E722E67E01A89 : begin ID22BB0550BCC1515614C8142FADDA171 = IDA65D1282C0B7B2A86436F0450F882A3 ;
end IDA65D1282C0B7B2A86436F0450F882A3 : begin if (I24C403550AE065D7D1B7266142886226 ) ID22BB0550BCC1515614C8142FADDA171
= IBE3FC19439FEC0073D66B4DAC2FECC32 ; end default : begin end endcase end  always @(posedge ICCFB0F435B37370076102F325BC08D20
or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin if (~I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin I37A362329A50BFF771D5547766A00B10
<= 1'b0; I2CA2FB392686EFC907D0D5C7FFF051AD <= 1'b0; IBE5A77ED6624B1E16464A1925007FB7C <= 1'b0; ID0A5ECECBEC8CE692F380DDF069E842F
<= 32'b0; I1877CB8174894BB7A9732E91A1794AAA <= 1'b0; I7E04E8229BE60B48AAE3E1EB6511163A <= IBE3FC19439FEC0073D66B4DAC2FECC32 ;
I612E93B17FEB6E7AE6FD9448B52CA816 <= 1'b0; I95FD0A1F8137860FD05FEA74508A613F <= 11'b0; I09934DCB789133B6EE69ED6ABA942F05
<= 1'b0; I8D181359467F27637239CDAEE8A2F45A <= 1'b0; end else begin I37A362329A50BFF771D5547766A00B10 <= (I2CA2FB392686EFC907D0D5C7FFF051AD
^ IBE5A77ED6624B1E16464A1925007FB7C ) ? 1'b1 : (I37A362329A50BFF771D5547766A00B10 & ~I5EA9375131D29CCE63A1B4FB334D5BBD );
I2CA2FB392686EFC907D0D5C7FFF051AD <= I1C0271AD5E8E9E9164909E468AD0B212 ; IBE5A77ED6624B1E16464A1925007FB7C <= I2CA2FB392686EFC907D0D5C7FFF051AD ;
I1877CB8174894BB7A9732E91A1794AAA <= 1'b0; I7E04E8229BE60B48AAE3E1EB6511163A <= ID22BB0550BCC1515614C8142FADDA171 ;
I09934DCB789133B6EE69ED6ABA942F05 <= 1'b0; case (I7E04E8229BE60B48AAE3E1EB6511163A ) IA7E2C061B23F9C2D79751962637FF9F8
: begin ID0A5ECECBEC8CE692F380DDF069E842F <= {(IBC983AF54FD90EA2AA9E3DD139A3B818 | {5'b0, IE46783A1FBEFC54C8AE5AC3DF183049F }),
24'b0}; I612E93B17FEB6E7AE6FD9448B52CA816 <= 1'b1; I09934DCB789133B6EE69ED6ABA942F05 <= 1'b1; end I0FBF38AB1DE3B938794F64EFEB6EEF04
: begin ID0A5ECECBEC8CE692F380DDF069E842F [31:8] <= {I3C7A9FA839F554D8898020C4831479E2 , I74A0936EE8FD1443A2C6745A4F3F6B5E ,
3'b111, 8'b0}; case (I691085C332A55972BA4126AE83875679 ) I1A3B3F253A4CAA84340E1092DB0AD78B : begin ID0A5ECECBEC8CE692F380DDF069E842F [7:0]
<= (I2CA2FB392686EFC907D0D5C7FFF051AD ) ? I476BD51644D400EA02C9B74EB861DDDC : I961C4AFB4B34DE00139652E84686874B ;
end I496D2BA2FDE6A39BB367B7EC043A5D8A : begin ID0A5ECECBEC8CE692F380DDF069E842F [7:0] <= (I2CA2FB392686EFC907D0D5C7FFF051AD )
? IDC0F38FB5CB3DE22405E2C1C80579AD8 : I508C4D4DDDB2A017FA853AA88EB418B2 ; end I0C9CD4F205090AE575352138FEB9E0B5
: begin ID0A5ECECBEC8CE692F380DDF069E842F [7:0] <= (I2CA2FB392686EFC907D0D5C7FFF051AD ) ? I64BD3AC45F8233E09BF36BB23F632819
: I4247280CBF50D75967C778AF3206D432 ; end I5898D0798C075683D57F7DA612ED3F03 : begin ID0A5ECECBEC8CE692F380DDF069E842F [7:0]
<= (I2CA2FB392686EFC907D0D5C7FFF051AD ) ? I68321D6CE308BEC2F016764C8A9FCEA8 : I72BD5161F8A297C6D1D0560048EA1612 ;
end default : begin ID0A5ECECBEC8CE692F380DDF069E842F [7:0] <= I961C4AFB4B34DE00139652E84686874B ; end endcase end
I2512657214BD8CD9D7C9E46341FB6960 : begin ID0A5ECECBEC8CE692F380DDF069E842F <= 32'b0; end IA4F9276F2E3EF93B14F2B0FF3B2DDE74
: begin I1877CB8174894BB7A9732E91A1794AAA <= 1'b1; end I3AEAA310DC2EB1E6D2E2AB4DD0417BA2 : begin I612E93B17FEB6E7AE6FD9448B52CA816
<= 1'b0; end I9CFCF3FC76F8BCD4AA7E722E67E01A89 : begin ID0A5ECECBEC8CE692F380DDF069E842F <= 32'b0; I8D181359467F27637239CDAEE8A2F45A
<= 1'b1; end IDA65D1282C0B7B2A86436F0450F882A3 : begin I8D181359467F27637239CDAEE8A2F45A <= I8D181359467F27637239CDAEE8A2F45A
& ~I24C403550AE065D7D1B7266142886226 ; end default : begin end endcase end end endmodule 
  module IE37A0AF0C4EF574205CEC4FFC0E18B72 #( parameter IAB32DAC10CBDBE04FD5EDBF7A576CAF9 = 512, I5F8A137EF3A5FDA6F2493F06E8FA441C
= 8 ) ( input wire ICCFB0F435B37370076102F325BC08D20 , input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire
IAE2A512A6B19FC0C3730E2011E6005C2 , input wire IB982FFD48AC89FC36697FE056A557C32 , input wire IBE1B10B19E9615FD92C8399CFD660D2E ,
input wire [I5F8A137EF3A5FDA6F2493F06E8FA441C - 1:0] I91C25096707DEBEF0FC17788A26B01A1 , input wire [I5F8A137EF3A5FDA6F2493F06E8FA441C
- 1:0] I6777AFB972CFFDA974EE962374CC84A0 , input wire [I5F8A137EF3A5FDA6F2493F06E8FA441C - 1:0] IA29FAC409EB1AFED4EA6D47BD6948E58 ,
input wire [I5F8A137EF3A5FDA6F2493F06E8FA441C - 1:0] I0B0360E6CCAB0F48EC1A783DD6B25856 , input wire [$clog2(IAB32DAC10CBDBE04FD5EDBF7A576CAF9
+ 1) - 1:0] I3FF97406B3ED373B267711109A980AF9 , output wire [I5F8A137EF3A5FDA6F2493F06E8FA441C - 1:0] I39B913343A3C8C7ED94053B14CAC4B0B ,
output wire [I5F8A137EF3A5FDA6F2493F06E8FA441C - 1:0] ID721B306FF47217933BAF6C84043D7D0 , output wire IA985CB046A7CFFDE37DDE98DA1CB21E0 ,
output wire I9F56096443CA90A430FDB4D329777AA2 , output wire [I5F8A137EF3A5FDA6F2493F06E8FA441C - 1:0] IB7E86A59807B16D5CCDC9D84A551E14D
);  localparam I9D9DF821BFE16A28B9DF536E518AB961 = 7; localparam I71E2CCCF89605682E005659BFB7C03FC = $clog2(IAB32DAC10CBDBE04FD5EDBF7A576CAF9
+ 1);  reg [I5F8A137EF3A5FDA6F2493F06E8FA441C - 1:0] IAAA9503DC311CD70C1EF204DB4F19CED ; reg [I5F8A137EF3A5FDA6F2493F06E8FA441C
- 1:0] I31B24A0AE0FE318B06D6CB78032BDA46 ; reg I5CA274DA39A18C8F0BC2765A88594483 ; reg IA5D44BAB064B6DE388B506B76B7F5E1E ;
reg I72868482C0602ADF96E1640AFFF3A6F9 ; reg [I5F8A137EF3A5FDA6F2493F06E8FA441C - 1:0] I2E017D4FD4F96203BF74C0264C9F0352 ;
reg [I5F8A137EF3A5FDA6F2493F06E8FA441C - 1:0] I397896584BEC0D07B2708021C6D18692 ; reg [I5F8A137EF3A5FDA6F2493F06E8FA441C
- 1:0] I74D457515F508FEEEE0B484060E44CC4 ; reg [I5F8A137EF3A5FDA6F2493F06E8FA441C - 1:0] ICB9A20003273C74B5FC4F24E27BF0CA4 ;
reg [I5F8A137EF3A5FDA6F2493F06E8FA441C - 1:0] IF68B76EBDAD735F87E59242264B17A6B ; reg [I5F8A137EF3A5FDA6F2493F06E8FA441C
- 1:0] I26ECBEE523A574CADF8B0D4C5A1428F4 ; reg [I5F8A137EF3A5FDA6F2493F06E8FA441C - 1:0] IE8FC206FE9A6600857461B50905895F8 ;
reg [I71E2CCCF89605682E005659BFB7C03FC - 1:0] I8FD1BCF7BFA2E3E11393B854E1DB9C6F ; reg I898781AD66FCB0FA1FAF902E88271FB1 ;
wire [I5F8A137EF3A5FDA6F2493F06E8FA441C - 1:0] I10EDC2BC5CA630453290335BC0902655 ; wire [I5F8A137EF3A5FDA6F2493F06E8FA441C
- 1:0] IF5F76BF56E7821B2B0BCC1FA7DA7C00F ; genvar I24501E622BFA6932719D2F78F75F6270 ;  assign I39B913343A3C8C7ED94053B14CAC4B0B
= I10EDC2BC5CA630453290335BC0902655 ; assign ID721B306FF47217933BAF6C84043D7D0 = I31B24A0AE0FE318B06D6CB78032BDA46 ;
assign IB7E86A59807B16D5CCDC9D84A551E14D = I2E017D4FD4F96203BF74C0264C9F0352 ; assign IA985CB046A7CFFDE37DDE98DA1CB21E0
= I5CA274DA39A18C8F0BC2765A88594483 ; assign I9F56096443CA90A430FDB4D329777AA2 = I72868482C0602ADF96E1640AFFF3A6F9 ;
 assign I10EDC2BC5CA630453290335BC0902655 = I26ECBEE523A574CADF8B0D4C5A1428F4 & ~IE8FC206FE9A6600857461B50905895F8 ;
 generate    for (I24501E622BFA6932719D2F78F75F6270 = 0; I24501E622BFA6932719D2F78F75F6270 < I5F8A137EF3A5FDA6F2493F06E8FA441C ;
I24501E622BFA6932719D2F78F75F6270 = I24501E622BFA6932719D2F78F75F6270 + 1) if (I24501E622BFA6932719D2F78F75F6270
== 0) assign IF5F76BF56E7821B2B0BCC1FA7DA7C00F [I24501E622BFA6932719D2F78F75F6270 ] = IF68B76EBDAD735F87E59242264B17A6B [I24501E622BFA6932719D2F78F75F6270 ]
& ~IB982FFD48AC89FC36697FE056A557C32 & I898781AD66FCB0FA1FAF902E88271FB1 ; else assign IF5F76BF56E7821B2B0BCC1FA7DA7C00F [I24501E622BFA6932719D2F78F75F6270 ]
= IF68B76EBDAD735F87E59242264B17A6B [I24501E622BFA6932719D2F78F75F6270 ] & ~(|IF68B76EBDAD735F87E59242264B17A6B [I24501E622BFA6932719D2F78F75F6270
- 1:0]) & ~IB982FFD48AC89FC36697FE056A557C32 & I898781AD66FCB0FA1FAF902E88271FB1 ; endgenerate  always @(posedge
ICCFB0F435B37370076102F325BC08D20 or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin if (~I9ED2A9117D3AEAF54CBA7AD69083BCB7 )
begin IAAA9503DC311CD70C1EF204DB4F19CED <= {I5F8A137EF3A5FDA6F2493F06E8FA441C {1'b0}}; I31B24A0AE0FE318B06D6CB78032BDA46
<= {I5F8A137EF3A5FDA6F2493F06E8FA441C {1'b0}}; I5CA274DA39A18C8F0BC2765A88594483 <= 1'b0; IA5D44BAB064B6DE388B506B76B7F5E1E
<= 1'b0; I72868482C0602ADF96E1640AFFF3A6F9 <= 1'b0; I2E017D4FD4F96203BF74C0264C9F0352 <= {I5F8A137EF3A5FDA6F2493F06E8FA441C {1'b0}};
I397896584BEC0D07B2708021C6D18692 <= {I5F8A137EF3A5FDA6F2493F06E8FA441C {1'b0}}; I74D457515F508FEEEE0B484060E44CC4
<= {I5F8A137EF3A5FDA6F2493F06E8FA441C {1'b0}}; ICB9A20003273C74B5FC4F24E27BF0CA4 <= {I5F8A137EF3A5FDA6F2493F06E8FA441C {1'b0}};
IF68B76EBDAD735F87E59242264B17A6B <= {I5F8A137EF3A5FDA6F2493F06E8FA441C {1'b0}}; I26ECBEE523A574CADF8B0D4C5A1428F4
<= {I5F8A137EF3A5FDA6F2493F06E8FA441C {1'b0}}; IE8FC206FE9A6600857461B50905895F8 <= {I5F8A137EF3A5FDA6F2493F06E8FA441C {1'b0}};
I8FD1BCF7BFA2E3E11393B854E1DB9C6F <= {I71E2CCCF89605682E005659BFB7C03FC {1'b0}}; I898781AD66FCB0FA1FAF902E88271FB1
<= 1'b0; end else begin IAAA9503DC311CD70C1EF204DB4F19CED <= IF5F76BF56E7821B2B0BCC1FA7DA7C00F ; I5CA274DA39A18C8F0BC2765A88594483
<= ~IAE2A512A6B19FC0C3730E2011E6005C2 & ~I5CA274DA39A18C8F0BC2765A88594483 & ~IA5D44BAB064B6DE388B506B76B7F5E1E
& ~(|I31B24A0AE0FE318B06D6CB78032BDA46 ); IA5D44BAB064B6DE388B506B76B7F5E1E <= I5CA274DA39A18C8F0BC2765A88594483
| (IA5D44BAB064B6DE388B506B76B7F5E1E & ~IBE1B10B19E9615FD92C8399CFD660D2E ); I72868482C0602ADF96E1640AFFF3A6F9 <=
|I10EDC2BC5CA630453290335BC0902655 ; I2E017D4FD4F96203BF74C0264C9F0352 <= IAAA9503DC311CD70C1EF204DB4F19CED ; I397896584BEC0D07B2708021C6D18692
<= I6777AFB972CFFDA974EE962374CC84A0 ; I74D457515F508FEEEE0B484060E44CC4 <= I31B24A0AE0FE318B06D6CB78032BDA46 &
IA29FAC409EB1AFED4EA6D47BD6948E58 ; ICB9A20003273C74B5FC4F24E27BF0CA4 <= I91C25096707DEBEF0FC17788A26B01A1 ; IF68B76EBDAD735F87E59242264B17A6B
<= ICB9A20003273C74B5FC4F24E27BF0CA4 & ~I26ECBEE523A574CADF8B0D4C5A1428F4 ; I26ECBEE523A574CADF8B0D4C5A1428F4 <=
IF5F76BF56E7821B2B0BCC1FA7DA7C00F | (I26ECBEE523A574CADF8B0D4C5A1428F4 & ~I74D457515F508FEEEE0B484060E44CC4 & ~I397896584BEC0D07B2708021C6D18692 );
IE8FC206FE9A6600857461B50905895F8 <= I26ECBEE523A574CADF8B0D4C5A1428F4 ; I8FD1BCF7BFA2E3E11393B854E1DB9C6F <= I3FF97406B3ED373B267711109A980AF9 ;
 I898781AD66FCB0FA1FAF902E88271FB1 <= (I8FD1BCF7BFA2E3E11393B854E1DB9C6F > I9D9DF821BFE16A28B9DF536E518AB961 ) ?
1'b1 : 1'b0; if (IBE1B10B19E9615FD92C8399CFD660D2E ) I31B24A0AE0FE318B06D6CB78032BDA46 <= I0B0360E6CCAB0F48EC1A783DD6B25856 ;
else I31B24A0AE0FE318B06D6CB78032BDA46 <= I31B24A0AE0FE318B06D6CB78032BDA46 & ~I74D457515F508FEEEE0B484060E44CC4
& ~I397896584BEC0D07B2708021C6D18692 ; end end endmodule
 module IFF5E0986AB6F727F3EEDED75702CE45A #( parameter IAB32DAC10CBDBE04FD5EDBF7A576CAF9 = 512, parameter I5F8A137EF3A5FDA6F2493F06E8FA441C
= 8, parameter I66C185998F46A7148163982E39BCD296 = "ecp3" ) ( input wire ICCFB0F435B37370076102F325BC08D20 , input
wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire [$clog2(IAB32DAC10CBDBE04FD5EDBF7A576CAF9 + 1) - 1:0] I3FF97406B3ED373B267711109A980AF9 ,
input wire [I5F8A137EF3A5FDA6F2493F06E8FA441C - 1:0] I91C25096707DEBEF0FC17788A26B01A1 , input wire [I5F8A137EF3A5FDA6F2493F06E8FA441C
- 1:0] I6777AFB972CFFDA974EE962374CC84A0 , input wire [I5F8A137EF3A5FDA6F2493F06E8FA441C - 1:0] IA29FAC409EB1AFED4EA6D47BD6948E58 ,
output wire [I5F8A137EF3A5FDA6F2493F06E8FA441C - 1:0] I39B913343A3C8C7ED94053B14CAC4B0B , output wire [I5F8A137EF3A5FDA6F2493F06E8FA441C
- 1:0] ID721B306FF47217933BAF6C84043D7D0 );  wire IB9E48499F019496BF412340B127E1839 ; wire IE78549D1E654EB948529EAED65694232 ;
wire [I5F8A137EF3A5FDA6F2493F06E8FA441C -1:0] I20ADF3B6DAF81414767B787F3D3ECD7C ; wire I92BBE8F1DA3A7479A827A07ADAD790B0 ;
wire I57B0F0FAE1ED417C46C84E0BF5BBB77B ; wire [I5F8A137EF3A5FDA6F2493F06E8FA441C -1:0] IEAD6835430C7C3605C25347A4056A838 ;
wire IF04BEDCC6C3F0AE64FE5531D24835A27 ;  IE37A0AF0C4EF574205CEC4FFC0E18B72 #( .IAB32DAC10CBDBE04FD5EDBF7A576CAF9
(IAB32DAC10CBDBE04FD5EDBF7A576CAF9 ), .I5F8A137EF3A5FDA6F2493F06E8FA441C (I5F8A137EF3A5FDA6F2493F06E8FA441C ) )
IB420C4D1279F971E867FA537CA4D6E82 ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .IAE2A512A6B19FC0C3730E2011E6005C2 (I92BBE8F1DA3A7479A827A07ADAD790B0 ), .IB982FFD48AC89FC36697FE056A557C32
(I57B0F0FAE1ED417C46C84E0BF5BBB77B ), .IBE1B10B19E9615FD92C8399CFD660D2E (IF04BEDCC6C3F0AE64FE5531D24835A27 ), .I91C25096707DEBEF0FC17788A26B01A1
(I91C25096707DEBEF0FC17788A26B01A1 ), .I6777AFB972CFFDA974EE962374CC84A0 (I6777AFB972CFFDA974EE962374CC84A0 ), .IA29FAC409EB1AFED4EA6D47BD6948E58
(IA29FAC409EB1AFED4EA6D47BD6948E58 ), .I0B0360E6CCAB0F48EC1A783DD6B25856 (IEAD6835430C7C3605C25347A4056A838 ), .I3FF97406B3ED373B267711109A980AF9
(I3FF97406B3ED373B267711109A980AF9 ), .I39B913343A3C8C7ED94053B14CAC4B0B (I39B913343A3C8C7ED94053B14CAC4B0B ), .ID721B306FF47217933BAF6C84043D7D0
(ID721B306FF47217933BAF6C84043D7D0 ), .IA985CB046A7CFFDE37DDE98DA1CB21E0 (IB9E48499F019496BF412340B127E1839 ), .I9F56096443CA90A430FDB4D329777AA2
(IE78549D1E654EB948529EAED65694232 ), .IB7E86A59807B16D5CCDC9D84A551E14D (I20ADF3B6DAF81414767B787F3D3ECD7C ) );
IF4FD65273243DC47A72869EEEA639DCD #( .I7292F55C07BFD7FB8A60D29FFC186275 (I5F8A137EF3A5FDA6F2493F06E8FA441C ), .IB71844FFA3AB85FEF45EAB4D35395752
(I5F8A137EF3A5FDA6F2493F06E8FA441C ), .I66C185998F46A7148163982E39BCD296 (I66C185998F46A7148163982E39BCD296 ) )
I65EC869BD2E9A693496F1F2E16A7ABA9 ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .IC79EC9A9F373F4B71374BDF6EDD31DE6 (1'b0), .I48D61F5A0B5732A58912433B42CD9D0C
(IB9E48499F019496BF412340B127E1839 ), .I04BC24D2B6403E54A64DE9E6C9ABAA2B (I20ADF3B6DAF81414767B787F3D3ECD7C ), .IE315CDCA06C9620D5C0AB966E553F0C3
(IE78549D1E654EB948529EAED65694232 ), .I11CEFC90537A67CD1FF01400245362F2 (), .ID7FCE45A65ADDB17F91F73A1B506BB5B
(), .I125028C7446331521D0434C10E8B0007 (IEAD6835430C7C3605C25347A4056A838 ), .I8BB939FF2AFDE7B2A1E480DCB61CE354
(I92BBE8F1DA3A7479A827A07ADAD790B0 ), .I41C63F948E534C7ED9F2471A44C922B2 (), .I585F74DE05DD9C1C7070D6B4F6E181C2
(IF04BEDCC6C3F0AE64FE5531D24835A27 ), .I705C64753A50CDA034B5ACB332D71768 (), .I233E0C0C8E5150F0CD8258F276D93942
(), .IBE0D6810EBD63B5C428623C578CF6D3A (I57B0F0FAE1ED417C46C84E0BF5BBB77B ), .I115E90220158F08B0465E99D7F2561D3
() ); endmodule
 module IB692DAE41499E4B01D446B8B28C804EB #( parameter I8F2F3EE9FE4B702742B51120C0EDA11A = 0, I73ABD5619A9FB885445AC1E288EAF7F8
= 0, I28B2C4B454208AC784C97EA8274B9503 = 1, ID538F704AA7B227247264F05C613DABA = 0 ) ( input wire ICCFB0F435B37370076102F325BC08D20 ,
input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire [7:0] I3C7A9FA839F554D8898020C4831479E2 , input wire [4:0]
I74A0936EE8FD1443A2C6745A4F3F6B5E , input wire [31:0] I1C0271AD5E8E9E9164909E468AD0B212 , input wire [11:0] I3D49ADB3C231E0C52B4EE7C42AB0DF8B ,
input wire [3:0] IE789C637CC57CC8ECB73F88C9790C5E4 , input wire [31:0] I3C3096B9DAB1C65EA381C7E05B767FB3 , input
wire I684F27663FD8A3EFB4B2BC8B42792CD0 , input wire I7378609E0B803011E82F6C6ABE861625 , input wire I56148DDDF284443347FFCF4F9C3BE61A ,
input wire I24C403550AE065D7D1B7266142886226 , output wire [31:0] IB808853736ABE6034DB8E375F1F00E89 , output wire
[31:0] IFE4A8CBA73734C6F0F0A078027E053D4 , output wire ID7A2A8B1E9D92B60194D5FAFAAB15208 , output wire IF274FAF97F5BACD693913BB418717A9D ,
output wire ID95C13E7EE1CFE6A8743FF9E62C25873 , output wire [10:0] IC58E411F24D810EF60A7B8638ABCC0BB , output wire
I89CFFA73C7546481B72B0FB06D799AEE , output wire I270ED686C2EF2C1C8B5B55EC4A5AAE84 ); `include "pcisig_constants.v"
function automatic [7:0] I19B1AF0FE0B2BA44377813F5D2133538 (input [7:0] IA0D1DB4FFBE8A7CF1A8A586BA8A56E12 ); begin
I19B1AF0FE0B2BA44377813F5D2133538 = {IA0D1DB4FFBE8A7CF1A8A586BA8A56E12 [7] & ~(|IA0D1DB4FFBE8A7CF1A8A586BA8A56E12 [6:0]),
IA0D1DB4FFBE8A7CF1A8A586BA8A56E12 [6] & ~(|IA0D1DB4FFBE8A7CF1A8A586BA8A56E12 [5:0]), IA0D1DB4FFBE8A7CF1A8A586BA8A56E12 [5]
& ~(|IA0D1DB4FFBE8A7CF1A8A586BA8A56E12 [4:0]), IA0D1DB4FFBE8A7CF1A8A586BA8A56E12 [4] & ~(|IA0D1DB4FFBE8A7CF1A8A586BA8A56E12 [3:0]),
IA0D1DB4FFBE8A7CF1A8A586BA8A56E12 [3] & ~(|IA0D1DB4FFBE8A7CF1A8A586BA8A56E12 [2:0]), IA0D1DB4FFBE8A7CF1A8A586BA8A56E12 [2]
& ~(|IA0D1DB4FFBE8A7CF1A8A586BA8A56E12 [1:0]), IA0D1DB4FFBE8A7CF1A8A586BA8A56E12 [1] & ~IA0D1DB4FFBE8A7CF1A8A586BA8A56E12 [0],
IA0D1DB4FFBE8A7CF1A8A586BA8A56E12 [0]}; end endfunction  reg [3:0] IF6762A005DECEE1D2D7F163C75BFEEC4 ; reg [31:0]
I0D2855032974DCC33735D9F8C9CAAA30 ; reg [31:0] IE2A4F3A7450FC95A7F9FF36380D08CEC ; reg [31:0] I3758FC83A1B5ACD9E6F20C2052725F78 ;
reg [4:0] I3D06B59E9F972357D2C9F413D0AD6BC8 ; reg [31:0] I2CA2FB392686EFC907D0D5C7FFF051AD ; reg [31:0] I349A82487A253B35E37EFDC7DAEF7F62 ;
reg [31:0] I454DE6E1D815566AC7AE0D064E785F96 ; reg [31:0] I543BA54CC3ABC74CF5E167DD24FC2851 ; reg [31:0] I2D40BAA904D8CD963B713EB1FBAC2D17 ;
reg I23ADFAC7E87DB224156796158F64B3F2 ; reg [3:0] IA41ECBBB6BB3AE10CC87C2948197DBF8 ; reg [3:0] IB9F6E6A6F23AFAFAC764389772A1B60D ;
reg [2:0] IF8856B01B16C2AAF77FFC519A21FACCC ; reg [4:0] I8E3E3A01C22724566C6D9D4F0D61A011 ; reg [7:0] I5443E4A5B263B816648B0A53C6158A99 ;
reg [31:0] I72E47AC634CDDC2338CBBD5642F81090 ; reg [31:0] I6ACE98A18452CD5394A3C8B4583C68B9 ; reg [31:0] IE10C2D271B10BCBDD51ACC08364CF5A2 ;
reg [31:0] I696440664361E19595FC920398AFDC38 ; reg [15:0] I54914F2A3BF3DCF1F71C331952F7B6C0 ; reg [31:0] ID0A5ECECBEC8CE692F380DDF069E842F ;
reg I1877CB8174894BB7A9732E91A1794AAA ; reg I612E93B17FEB6E7AE6FD9448B52CA816 ; reg [10:0] I95FD0A1F8137860FD05FEA74508A613F ;
reg I09934DCB789133B6EE69ED6ABA942F05 ; reg I8D181359467F27637239CDAEE8A2F45A ; wire [31:0] I91047088394D6A4116575942899FC337 ;
wire [31:0] IBC9BBA91B18A09BDF37FAB697B1D125B ; wire [11:0] IDF2D2EFCFCAA060A180881D81395C002 ; wire IBD4351E5DD0E0A5E0B00AA0548196F09 ;
 localparam I65DDC49F11A5CEA91E63CED60C1D3A4A = 4'b0000, I647611C5549265C57828CEEDA18C31A9 = 4'b0001, ID0A1D3F69F0CE541B268BDF88CB8EC16
= 4'b0010, I3B3571D42B3E5DB00256EFEF03B0C9A1 = 4'b0011, IDA78053AE36FF6CFD201CDBEA506FA6F = 4'b0100, I540E4DFE1B15CB8C9E38CD199B3772B8
= 4'b0101, I5900903CDB155403F0AFD0EA873FED3B = 4'b0110, I3A013BF4B9D3A78D76EB9E243941F7A8 = 4'b0111, ID1DB35908E01690E4664B488CAFF89AE
= 4'b1000, I2DCDAE01131E1BC9349FC6E12C6A7B49 = 4'b1001, IC5EAA87AE409D7C8DBF971ECD27F0F48 = 4'b1010; localparam
[2:0] I2349891C690C1942F0AB29644BF3A949 = I73ABD5619A9FB885445AC1E288EAF7F8 ;  localparam [15:0] I0A12D06C0E7540345D5CFBCA668D8E45
= (I28B2C4B454208AC784C97EA8274B9503 > 16) ? 16'h008a : ((I28B2C4B454208AC784C97EA8274B9503 > 8) ? 16'h0088 : ((I28B2C4B454208AC784C97EA8274B9503
> 4) ? 16'h0086 : ((I28B2C4B454208AC784C97EA8274B9503 > 2) ? 16'h0084 : ((I28B2C4B454208AC784C97EA8274B9503 > 1)
? 16'h0082 : 16'h0080)))); localparam [31:0] I275DFC10FBB3E818C9C99DF4FF58164C = 32'hffff0000; localparam [31:0]
IB3B48366BD64A201301128D3C38A67E9 = 32'hff00ff00; localparam [31:0] I7402C4BC57ED69FBAECF82EF36182142 = 32'hf0f0f0f0;
localparam [31:0] IBB94BBEBA5FFE253FAECF658F4B53993 = 32'hcccccccc; localparam [31:0] I844463A9769B79933942580A194992D1
= 32'haaaaaaaa; localparam [31:0] I4CD0CE6E86D910B226DA70EB032DFC85 = 32'h55555555; localparam [31:0] I0FEAB7D3056FDE01396D69D7687C9DDB
= 32'h01010101; localparam [31:0] I15AC5D8E5AEEF46487350EEEA52D84AE = 32'h02020202; localparam [31:0] IF2EB38FF515658D58F564B69266D3C12
= 32'h04040404; localparam [31:0] I51F14E3CFED73228615FAE55DED33499 = 32'h08080808; localparam [31:0] I1FF060A34E9842AA554A3F6838FDECEF
= 32'h10101010; localparam [31:0] IF754C10545FBD28AF98C3E8DABE1625F = 32'h20202020; localparam [31:0] I996C241A0424B970A2D6C63C55615E7F
= 32'h40404040; localparam [31:0] I68AE95FD8EAA7E7FA01B800C88945BF5 = 32'h80808080; localparam [31:0] IF83F67C5A73A1BB7CF01F279B6F2C858
= 32'h11111111; localparam [31:0] I6501B441F3CCC90245533CC5EEDABC4D = 32'h22222222; localparam [31:0] IC5FC1A4F5407EC9E61EA193A2ABD065B
= 32'h44444444; localparam [31:0] I08AE85FA7B91C13FA36E8E7CC0D74E8E = 32'h88888888; localparam [31:0] I1319A9AA88F5409F43101FB338E31183
= 32'haaaaaaaa; localparam [15:0] I1314FF8642ED3882C856F80D07EFA905 = 16'h0080; localparam [15:0] ID7692E171623C59210D3CCFC10E1B208
= 16'hff8e; localparam [7:0] I6D17E9EDD00B4065D8E70000AC734145 = ID538F704AA7B227247264F05C613DABA ; localparam
[11:0] I4D1E7463132962B155070B6AB1A37C8F = I8F2F3EE9FE4B702742B51120C0EDA11A + 12'h000; localparam [11:0] I95B7675879933B29B289575BCCB50121
= (I1314FF8642ED3882C856F80D07EFA905 [7] == 1'b1) ? (I8F2F3EE9FE4B702742B51120C0EDA11A + 12'h008) : (I8F2F3EE9FE4B702742B51120C0EDA11A
+ 12'hffc); localparam [11:0] I5B35B9EB726C2B745F5F926AAE3EF6AD = I8F2F3EE9FE4B702742B51120C0EDA11A + 12'h004; localparam
[11:0] I48D66DC51DBC9EB60A39D68068788DB9 = (I1314FF8642ED3882C856F80D07EFA905 [7] == 1'b1) ? (I8F2F3EE9FE4B702742B51120C0EDA11A
+ 12'h00c) : (I8F2F3EE9FE4B702742B51120C0EDA11A + 12'h008);  assign IB808853736ABE6034DB8E375F1F00E89 = I7378609E0B803011E82F6C6ABE861625
? I72E47AC634CDDC2338CBBD5642F81090 : 32'b0; assign IFE4A8CBA73734C6F0F0A078027E053D4 = ID0A5ECECBEC8CE692F380DDF069E842F ;
assign ID7A2A8B1E9D92B60194D5FAFAAB15208 = I1877CB8174894BB7A9732E91A1794AAA ; assign IF274FAF97F5BACD693913BB418717A9D
= I612E93B17FEB6E7AE6FD9448B52CA816 ; assign ID95C13E7EE1CFE6A8743FF9E62C25873 = IBD4351E5DD0E0A5E0B00AA0548196F09 ;
assign IC58E411F24D810EF60A7B8638ABCC0BB = I95FD0A1F8137860FD05FEA74508A613F ; assign I89CFFA73C7546481B72B0FB06D799AEE
= I09934DCB789133B6EE69ED6ABA942F05 ; assign I270ED686C2EF2C1C8B5B55EC4A5AAE84 = I8D181359467F27637239CDAEE8A2F45A ;
 assign I91047088394D6A4116575942899FC337 = I543BA54CC3ABC74CF5E167DD24FC2851 & ~I2D40BAA904D8CD963B713EB1FBAC2D17 ;
assign IBC9BBA91B18A09BDF37FAB697B1D125B = (I696440664361E19595FC920398AFDC38 & {{27{1'b1}}, I5443E4A5B263B816648B0A53C6158A99 [4:0]})
| ({27'b0, (~I5443E4A5B263B816648B0A53C6158A99 [4:0] & I8E3E3A01C22724566C6D9D4F0D61A011 )}); assign IDF2D2EFCFCAA060A180881D81395C002
= I3D49ADB3C231E0C52B4EE7C42AB0DF8B & 12'hffc; assign IBD4351E5DD0E0A5E0B00AA0548196F09 = (IA41ECBBB6BB3AE10CC87C2948197DBF8
== I3B3571D42B3E5DB00256EFEF03B0C9A1 ) ? 1'b1 : 1'b0;  always @(I2CA2FB392686EFC907D0D5C7FFF051AD or I454DE6E1D815566AC7AE0D064E785F96
or I23ADFAC7E87DB224156796158F64B3F2 or IA41ECBBB6BB3AE10CC87C2948197DBF8 or I6ACE98A18452CD5394A3C8B4583C68B9 or
I56148DDDF284443347FFCF4F9C3BE61A or I24C403550AE065D7D1B7266142886226 ) begin IB9F6E6A6F23AFAFAC764389772A1B60D
= IA41ECBBB6BB3AE10CC87C2948197DBF8 ; case (IA41ECBBB6BB3AE10CC87C2948197DBF8 ) I65DDC49F11A5CEA91E63CED60C1D3A4A
: begin if (I23ADFAC7E87DB224156796158F64B3F2 & (|I2CA2FB392686EFC907D0D5C7FFF051AD )) IB9F6E6A6F23AFAFAC764389772A1B60D
= I647611C5549265C57828CEEDA18C31A9 ; end I647611C5549265C57828CEEDA18C31A9 : begin IB9F6E6A6F23AFAFAC764389772A1B60D
= ID0A1D3F69F0CE541B268BDF88CB8EC16 ; end ID0A1D3F69F0CE541B268BDF88CB8EC16 : begin if (I454DE6E1D815566AC7AE0D064E785F96 )
IB9F6E6A6F23AFAFAC764389772A1B60D = I3B3571D42B3E5DB00256EFEF03B0C9A1 ; else IB9F6E6A6F23AFAFAC764389772A1B60D =
I65DDC49F11A5CEA91E63CED60C1D3A4A ; end I3B3571D42B3E5DB00256EFEF03B0C9A1 : begin if (I56148DDDF284443347FFCF4F9C3BE61A )
IB9F6E6A6F23AFAFAC764389772A1B60D = IDA78053AE36FF6CFD201CDBEA506FA6F ; end IDA78053AE36FF6CFD201CDBEA506FA6F :
begin IB9F6E6A6F23AFAFAC764389772A1B60D = I540E4DFE1B15CB8C9E38CD199B3772B8 ; end I540E4DFE1B15CB8C9E38CD199B3772B8
: begin IB9F6E6A6F23AFAFAC764389772A1B60D = I5900903CDB155403F0AFD0EA873FED3B ; end I5900903CDB155403F0AFD0EA873FED3B
: begin IB9F6E6A6F23AFAFAC764389772A1B60D = I3A013BF4B9D3A78D76EB9E243941F7A8 ; end I3A013BF4B9D3A78D76EB9E243941F7A8
: begin if (I6ACE98A18452CD5394A3C8B4583C68B9 ) IB9F6E6A6F23AFAFAC764389772A1B60D = ID1DB35908E01690E4664B488CAFF89AE ;
else IB9F6E6A6F23AFAFAC764389772A1B60D = I2DCDAE01131E1BC9349FC6E12C6A7B49 ; end ID1DB35908E01690E4664B488CAFF89AE
: begin IB9F6E6A6F23AFAFAC764389772A1B60D = I2DCDAE01131E1BC9349FC6E12C6A7B49 ; end I2DCDAE01131E1BC9349FC6E12C6A7B49
: begin IB9F6E6A6F23AFAFAC764389772A1B60D = IC5EAA87AE409D7C8DBF971ECD27F0F48 ; end IC5EAA87AE409D7C8DBF971ECD27F0F48
: begin if (I24C403550AE065D7D1B7266142886226 ) IB9F6E6A6F23AFAFAC764389772A1B60D = ID0A1D3F69F0CE541B268BDF88CB8EC16 ;
end default : begin end endcase end  always @(IDF2D2EFCFCAA060A180881D81395C002 or I7378609E0B803011E82F6C6ABE861625 )
begin  if (I7378609E0B803011E82F6C6ABE861625 ) case (IDF2D2EFCFCAA060A180881D81395C002 ) I5B35B9EB726C2B745F5F926AAE3EF6AD
: I72E47AC634CDDC2338CBBD5642F81090 = IE10C2D271B10BCBDD51ACC08364CF5A2 ; I95B7675879933B29B289575BCCB50121 : I72E47AC634CDDC2338CBBD5642F81090
= (I1314FF8642ED3882C856F80D07EFA905 [7] == 1'b1) ? I6ACE98A18452CD5394A3C8B4583C68B9 : 32'b0; I48D66DC51DBC9EB60A39D68068788DB9
: I72E47AC634CDDC2338CBBD5642F81090 = I696440664361E19595FC920398AFDC38 ; I4D1E7463132962B155070B6AB1A37C8F : I72E47AC634CDDC2338CBBD5642F81090
= {(I54914F2A3BF3DCF1F71C331952F7B6C0 | I0A12D06C0E7540345D5CFBCA668D8E45 ), I6D17E9EDD00B4065D8E70000AC734145 ,
I92BEFE7DA8E3713D40B466EEDA052B30 }; default : I72E47AC634CDDC2338CBBD5642F81090 = 32'b0; endcase else I72E47AC634CDDC2338CBBD5642F81090
= 32'b0; end  always @(posedge ICCFB0F435B37370076102F325BC08D20 or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 )
begin if (~I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin IF6762A005DECEE1D2D7F163C75BFEEC4 <= 4'b0; I0D2855032974DCC33735D9F8C9CAAA30
<= 32'b0; IE2A4F3A7450FC95A7F9FF36380D08CEC <= 32'b0; I3758FC83A1B5ACD9E6F20C2052725F78 <= 32'b0; I3D06B59E9F972357D2C9F413D0AD6BC8
<= 5'b0; I2CA2FB392686EFC907D0D5C7FFF051AD <= 32'b0; I349A82487A253B35E37EFDC7DAEF7F62 <= 32'b0; I454DE6E1D815566AC7AE0D064E785F96
<= 32'b0; I543BA54CC3ABC74CF5E167DD24FC2851 <= 32'b0; I2D40BAA904D8CD963B713EB1FBAC2D17 <= 32'b0; I23ADFAC7E87DB224156796158F64B3F2
<= 1'b0; IA41ECBBB6BB3AE10CC87C2948197DBF8 <= 4'b0; IF8856B01B16C2AAF77FFC519A21FACCC <= 3'b0; I8E3E3A01C22724566C6D9D4F0D61A011
<= 5'b0; I5443E4A5B263B816648B0A53C6158A99 <= 5'b0; I6ACE98A18452CD5394A3C8B4583C68B9 <= 32'b0; IE10C2D271B10BCBDD51ACC08364CF5A2
<= 32'b0; I54914F2A3BF3DCF1F71C331952F7B6C0 <= I1314FF8642ED3882C856F80D07EFA905 & ID7692E171623C59210D3CCFC10E1B208 ;
I696440664361E19595FC920398AFDC38 <= 32'b0; ID0A5ECECBEC8CE692F380DDF069E842F <= 32'b0; I1877CB8174894BB7A9732E91A1794AAA
<= 1'b0; I612E93B17FEB6E7AE6FD9448B52CA816 <= 1'b0; I95FD0A1F8137860FD05FEA74508A613F <= 11'b0; I09934DCB789133B6EE69ED6ABA942F05
<= 1'b0; I8D181359467F27637239CDAEE8A2F45A <= 1'b0; end else begin    IF6762A005DECEE1D2D7F163C75BFEEC4 <= {|I454DE6E1D815566AC7AE0D064E785F96 [31:24],
|I454DE6E1D815566AC7AE0D064E785F96 [23:16], |I454DE6E1D815566AC7AE0D064E785F96 [15:8], |I454DE6E1D815566AC7AE0D064E785F96 [7:0]};
I0D2855032974DCC33735D9F8C9CAAA30 <= {I19B1AF0FE0B2BA44377813F5D2133538 (I454DE6E1D815566AC7AE0D064E785F96 [31:24]),
I19B1AF0FE0B2BA44377813F5D2133538 (I454DE6E1D815566AC7AE0D064E785F96 [23:16]), I19B1AF0FE0B2BA44377813F5D2133538 (I454DE6E1D815566AC7AE0D064E785F96 [15:8]),
I19B1AF0FE0B2BA44377813F5D2133538 (I454DE6E1D815566AC7AE0D064E785F96 [7:0])}; IE2A4F3A7450FC95A7F9FF36380D08CEC
<= {((|IF6762A005DECEE1D2D7F163C75BFEEC4 [2:0]) ? 8'b00 : I0D2855032974DCC33735D9F8C9CAAA30 [31:24]), ((|IF6762A005DECEE1D2D7F163C75BFEEC4 [1:0])
? 8'b00 : I0D2855032974DCC33735D9F8C9CAAA30 [23:16]), ((IF6762A005DECEE1D2D7F163C75BFEEC4 [0]) ? 8'b00 : I0D2855032974DCC33735D9F8C9CAAA30 [15:8]),
I0D2855032974DCC33735D9F8C9CAAA30 [7:0]}; I3758FC83A1B5ACD9E6F20C2052725F78 <= (IB9F6E6A6F23AFAFAC764389772A1B60D
== I2DCDAE01131E1BC9349FC6E12C6A7B49 ) ? IE2A4F3A7450FC95A7F9FF36380D08CEC : 32'b0; I2CA2FB392686EFC907D0D5C7FFF051AD
<= I91047088394D6A4116575942899FC337 | (I2CA2FB392686EFC907D0D5C7FFF051AD & ~I3758FC83A1B5ACD9E6F20C2052725F78 );
I349A82487A253B35E37EFDC7DAEF7F62 <= I1C0271AD5E8E9E9164909E468AD0B212 ; I454DE6E1D815566AC7AE0D064E785F96 <= (IA41ECBBB6BB3AE10CC87C2948197DBF8
== I647611C5549265C57828CEEDA18C31A9 ) ? I2CA2FB392686EFC907D0D5C7FFF051AD : (I454DE6E1D815566AC7AE0D064E785F96
& ~I3758FC83A1B5ACD9E6F20C2052725F78 ); I2D40BAA904D8CD963B713EB1FBAC2D17 <= I543BA54CC3ABC74CF5E167DD24FC2851 ;
I23ADFAC7E87DB224156796158F64B3F2 <= I54914F2A3BF3DCF1F71C331952F7B6C0 [0]; IA41ECBBB6BB3AE10CC87C2948197DBF8 <=
IB9F6E6A6F23AFAFAC764389772A1B60D ; IF8856B01B16C2AAF77FFC519A21FACCC <= I54914F2A3BF3DCF1F71C331952F7B6C0 [6:4];
I8E3E3A01C22724566C6D9D4F0D61A011 [4] <= |(IE2A4F3A7450FC95A7F9FF36380D08CEC & I275DFC10FBB3E818C9C99DF4FF58164C );
I8E3E3A01C22724566C6D9D4F0D61A011 [3] <= |(IE2A4F3A7450FC95A7F9FF36380D08CEC & IB3B48366BD64A201301128D3C38A67E9 );
I8E3E3A01C22724566C6D9D4F0D61A011 [2] <= |(IE2A4F3A7450FC95A7F9FF36380D08CEC & I7402C4BC57ED69FBAECF82EF36182142 );
I8E3E3A01C22724566C6D9D4F0D61A011 [1] <= |(IE2A4F3A7450FC95A7F9FF36380D08CEC & IBB94BBEBA5FFE253FAECF658F4B53993 );
I8E3E3A01C22724566C6D9D4F0D61A011 [0] <= |(IE2A4F3A7450FC95A7F9FF36380D08CEC & I844463A9769B79933942580A194992D1 );
 case (IF8856B01B16C2AAF77FFC519A21FACCC ) 3'b000 : begin I543BA54CC3ABC74CF5E167DD24FC2851 <= {31'b0, |I349A82487A253B35E37EFDC7DAEF7F62 };
I5443E4A5B263B816648B0A53C6158A99 <= 8'hff; end 3'b001 : begin I543BA54CC3ABC74CF5E167DD24FC2851 <= {30'b0, |(I349A82487A253B35E37EFDC7DAEF7F62
& I1319A9AA88F5409F43101FB338E31183 ), |(I349A82487A253B35E37EFDC7DAEF7F62 & I4CD0CE6E86D910B226DA70EB032DFC85 )};
I5443E4A5B263B816648B0A53C6158A99 <= 8'hfe; end 3'b010 : begin I543BA54CC3ABC74CF5E167DD24FC2851 <= {28'b0, |(I349A82487A253B35E37EFDC7DAEF7F62
& I08AE85FA7B91C13FA36E8E7CC0D74E8E ), |(I349A82487A253B35E37EFDC7DAEF7F62 & IC5FC1A4F5407EC9E61EA193A2ABD065B ),
|(I349A82487A253B35E37EFDC7DAEF7F62 & I6501B441F3CCC90245533CC5EEDABC4D ), |(I349A82487A253B35E37EFDC7DAEF7F62 &
IF83F67C5A73A1BB7CF01F279B6F2C858 )}; I5443E4A5B263B816648B0A53C6158A99 <= 8'hfc; end 3'b011 : begin I543BA54CC3ABC74CF5E167DD24FC2851
<= {24'b0, |(I349A82487A253B35E37EFDC7DAEF7F62 & I68AE95FD8EAA7E7FA01B800C88945BF5 ), |(I349A82487A253B35E37EFDC7DAEF7F62
& I996C241A0424B970A2D6C63C55615E7F ), |(I349A82487A253B35E37EFDC7DAEF7F62 & IF754C10545FBD28AF98C3E8DABE1625F ),
|(I349A82487A253B35E37EFDC7DAEF7F62 & I1FF060A34E9842AA554A3F6838FDECEF ), |(I349A82487A253B35E37EFDC7DAEF7F62 &
I51F14E3CFED73228615FAE55DED33499 ), |(I349A82487A253B35E37EFDC7DAEF7F62 & IF2EB38FF515658D58F564B69266D3C12 ),
|(I349A82487A253B35E37EFDC7DAEF7F62 & I15AC5D8E5AEEF46487350EEEA52D84AE ), |(I349A82487A253B35E37EFDC7DAEF7F62 &
I0FEAB7D3056FDE01396D69D7687C9DDB )}; I5443E4A5B263B816648B0A53C6158A99 <= 8'hf8; end 3'b100 : begin I543BA54CC3ABC74CF5E167DD24FC2851
<= {16'b0, (I349A82487A253B35E37EFDC7DAEF7F62 [31:16] | I349A82487A253B35E37EFDC7DAEF7F62 [15:0])}; I5443E4A5B263B816648B0A53C6158A99
<= 8'hf0; end default : begin I543BA54CC3ABC74CF5E167DD24FC2851 <= I349A82487A253B35E37EFDC7DAEF7F62 ; I5443E4A5B263B816648B0A53C6158A99
<= 8'he0; end endcase  case (IA41ECBBB6BB3AE10CC87C2948197DBF8 ) ID0A1D3F69F0CE541B268BDF88CB8EC16 : begin I95FD0A1F8137860FD05FEA74508A613F
<= 11'h001; end IDA78053AE36FF6CFD201CDBEA506FA6F : begin ID0A5ECECBEC8CE692F380DDF069E842F <= (I6ACE98A18452CD5394A3C8B4583C68B9 )
? {I2E664E814B6AA2CBCE57FBCE2A354435 , 16'b0, 8'h01} : {IEC10F95DD42CAF869EFB03BDF59BE8EB , 16'b0, 8'h01}; I612E93B17FEB6E7AE6FD9448B52CA816
<= 1'b1; I09934DCB789133B6EE69ED6ABA942F05 <= 1'b1; end I540E4DFE1B15CB8C9E38CD199B3772B8 : begin ID0A5ECECBEC8CE692F380DDF069E842F
<= {I3C7A9FA839F554D8898020C4831479E2 , I74A0936EE8FD1443A2C6745A4F3F6B5E , I2349891C690C1942F0AB29644BF3A949 ,
8'b0, 8'h03}; I09934DCB789133B6EE69ED6ABA942F05 <= 1'b0; end I5900903CDB155403F0AFD0EA873FED3B : ID0A5ECECBEC8CE692F380DDF069E842F
<= (I6ACE98A18452CD5394A3C8B4583C68B9 ) ? I6ACE98A18452CD5394A3C8B4583C68B9 : IE10C2D271B10BCBDD51ACC08364CF5A2 ;
I3A013BF4B9D3A78D76EB9E243941F7A8 : begin ID0A5ECECBEC8CE692F380DDF069E842F <= (I6ACE98A18452CD5394A3C8B4583C68B9 )
? IE10C2D271B10BCBDD51ACC08364CF5A2 : {IBC9BBA91B18A09BDF37FAB697B1D125B [7:0], IBC9BBA91B18A09BDF37FAB697B1D125B [15:8],
IBC9BBA91B18A09BDF37FAB697B1D125B [23:16], IBC9BBA91B18A09BDF37FAB697B1D125B [31:24]}; I1877CB8174894BB7A9732E91A1794AAA
<= (I6ACE98A18452CD5394A3C8B4583C68B9 ) ? 1'b0 : 1'b1; end ID1DB35908E01690E4664B488CAFF89AE : begin ID0A5ECECBEC8CE692F380DDF069E842F
<= {IBC9BBA91B18A09BDF37FAB697B1D125B [7:0], IBC9BBA91B18A09BDF37FAB697B1D125B [15:8], IBC9BBA91B18A09BDF37FAB697B1D125B [23:16],
IBC9BBA91B18A09BDF37FAB697B1D125B [31:24]}; I1877CB8174894BB7A9732E91A1794AAA <= 1'b1; end I2DCDAE01131E1BC9349FC6E12C6A7B49
: begin ID0A5ECECBEC8CE692F380DDF069E842F <= 32'b0; I1877CB8174894BB7A9732E91A1794AAA <= 1'b0; I612E93B17FEB6E7AE6FD9448B52CA816
<= 1'b0; I8D181359467F27637239CDAEE8A2F45A <= 1'b1; end IC5EAA87AE409D7C8DBF971ECD27F0F48 : begin I95FD0A1F8137860FD05FEA74508A613F
<= 11'b0; I8D181359467F27637239CDAEE8A2F45A <= I8D181359467F27637239CDAEE8A2F45A & ~I24C403550AE065D7D1B7266142886226 ;
end default : begin end endcase  if (I7378609E0B803011E82F6C6ABE861625 & I684F27663FD8A3EFB4B2BC8B42792CD0 ) begin
case (IDF2D2EFCFCAA060A180881D81395C002 ) I5B35B9EB726C2B745F5F926AAE3EF6AD : begin if (IE789C637CC57CC8ECB73F88C9790C5E4 [0])
IE10C2D271B10BCBDD51ACC08364CF5A2 [7:0] <= I3C3096B9DAB1C65EA381C7E05B767FB3 [7:0]; if (IE789C637CC57CC8ECB73F88C9790C5E4 [1])
IE10C2D271B10BCBDD51ACC08364CF5A2 [15:8] <= I3C3096B9DAB1C65EA381C7E05B767FB3 [15:8]; if (IE789C637CC57CC8ECB73F88C9790C5E4 [2])
IE10C2D271B10BCBDD51ACC08364CF5A2 [23:15] <= I3C3096B9DAB1C65EA381C7E05B767FB3 [23:15]; if (IE789C637CC57CC8ECB73F88C9790C5E4 [3])
IE10C2D271B10BCBDD51ACC08364CF5A2 [31:24] <= I3C3096B9DAB1C65EA381C7E05B767FB3 [31:24]; end I95B7675879933B29B289575BCCB50121
: begin if (I1314FF8642ED3882C856F80D07EFA905 [0] == 1'b1) begin if (IE789C637CC57CC8ECB73F88C9790C5E4 [0]) I6ACE98A18452CD5394A3C8B4583C68B9 [7:0]
<= I3C3096B9DAB1C65EA381C7E05B767FB3 [7:0]; if (IE789C637CC57CC8ECB73F88C9790C5E4 [1]) I6ACE98A18452CD5394A3C8B4583C68B9 [15:8]
<= I3C3096B9DAB1C65EA381C7E05B767FB3 [15:8]; if (IE789C637CC57CC8ECB73F88C9790C5E4 [2]) I6ACE98A18452CD5394A3C8B4583C68B9 [23:15]
<= I3C3096B9DAB1C65EA381C7E05B767FB3 [23:15]; if (IE789C637CC57CC8ECB73F88C9790C5E4 [3]) I6ACE98A18452CD5394A3C8B4583C68B9 [31:24]
<= I3C3096B9DAB1C65EA381C7E05B767FB3 [31:24]; end end I48D66DC51DBC9EB60A39D68068788DB9 : begin if (IE789C637CC57CC8ECB73F88C9790C5E4 [0])
I696440664361E19595FC920398AFDC38 [7:0] <= I3C3096B9DAB1C65EA381C7E05B767FB3 [7:0] & I5443E4A5B263B816648B0A53C6158A99 ;
if (IE789C637CC57CC8ECB73F88C9790C5E4 [1]) I696440664361E19595FC920398AFDC38 [15:8] <= I3C3096B9DAB1C65EA381C7E05B767FB3 [15:8];
if (IE789C637CC57CC8ECB73F88C9790C5E4 [2]) I696440664361E19595FC920398AFDC38 [23:15] <= I3C3096B9DAB1C65EA381C7E05B767FB3 [23:15];
if (IE789C637CC57CC8ECB73F88C9790C5E4 [3]) I696440664361E19595FC920398AFDC38 [31:24] <= I3C3096B9DAB1C65EA381C7E05B767FB3 [31:24];
end I4D1E7463132962B155070B6AB1A37C8F : begin if (IE789C637CC57CC8ECB73F88C9790C5E4 [2]) I54914F2A3BF3DCF1F71C331952F7B6C0 [7:0]
<= (I54914F2A3BF3DCF1F71C331952F7B6C0 [7:0] & ID7692E171623C59210D3CCFC10E1B208 [7:0]) | (I3C3096B9DAB1C65EA381C7E05B767FB3 [23:16]
& ~ID7692E171623C59210D3CCFC10E1B208 [7:0]); if (IE789C637CC57CC8ECB73F88C9790C5E4 [3]) I54914F2A3BF3DCF1F71C331952F7B6C0 [15:8]
<= (I54914F2A3BF3DCF1F71C331952F7B6C0 [15:8] & ID7692E171623C59210D3CCFC10E1B208 [15:8]) | (I3C3096B9DAB1C65EA381C7E05B767FB3 [31:24]
& ~ID7692E171623C59210D3CCFC10E1B208 [15:8]); end endcase end end end endmodule 
 module IF44E5E7AB65AFFA1AF3DA949DB91C839 #( parameter I8F2F3EE9FE4B702742B51120C0EDA11A = 0, ID538F704AA7B227247264F05C613DABA
= 0 ) ( input wire ICCFB0F435B37370076102F325BC08D20 , input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire
[11:0] I3D49ADB3C231E0C52B4EE7C42AB0DF8B , input wire [3:0] IE789C637CC57CC8ECB73F88C9790C5E4 , input wire [31:0]
I3C3096B9DAB1C65EA381C7E05B767FB3 , input wire I684F27663FD8A3EFB4B2BC8B42792CD0 , input wire I7378609E0B803011E82F6C6ABE861625 ,
output wire I31CF69FF368B36B4D6612DF16B3ABC6B , output wire I26F316E89E4B007444B724CD95758235 , output wire [31:0]
IB808853736ABE6034DB8E375F1F00E89 ); `include "pcisig_constants.v"
 reg I9B8138DCE156F7C31EB5914EF01F183C ; reg IFFD0BAB32DEE73305A584A062E784936 ; reg [31:0] I72E47AC634CDDC2338CBBD5642F81090 ;
reg [15:0] I9C49DC380ED90CDC0B86D16428C58A39 ; wire [11:0] I50BC02B32FFEA3FDDA09A1A76C72EDE6 ; wire [11:0] I23CD01FB20FA1C856A43C90DA2FE8B37 ;
wire [7:0] IB733A674E6EDACC67D7A142D9C749704 ; wire [11:0] IDF2D2EFCFCAA060A180881D81395C002 ;  localparam I14E299D2F1F5A86F6DF0D7820BB0365E
= I8F2F3EE9FE4B702742B51120C0EDA11A + 12'h004;  localparam IDD2F1F37B45AD83BB6A8FD6BED814957 = 2'b00;  assign I31CF69FF368B36B4D6612DF16B3ABC6B
= I9B8138DCE156F7C31EB5914EF01F183C ; assign I26F316E89E4B007444B724CD95758235 = IFFD0BAB32DEE73305A584A062E784936 ;
assign IB808853736ABE6034DB8E375F1F00E89 = I7378609E0B803011E82F6C6ABE861625 ? I72E47AC634CDDC2338CBBD5642F81090
: 32'b0;  assign IDF2D2EFCFCAA060A180881D81395C002 = I3D49ADB3C231E0C52B4EE7C42AB0DF8B & 12'hffc; generate assign
I50BC02B32FFEA3FDDA09A1A76C72EDE6 = I14E299D2F1F5A86F6DF0D7820BB0365E ; assign I23CD01FB20FA1C856A43C90DA2FE8B37
= I8F2F3EE9FE4B702742B51120C0EDA11A ; assign IB733A674E6EDACC67D7A142D9C749704 = ID538F704AA7B227247264F05C613DABA ;
endgenerate  always @(IDF2D2EFCFCAA060A180881D81395C002 or I9C49DC380ED90CDC0B86D16428C58A39 or I7378609E0B803011E82F6C6ABE861625 )
begin if (I7378609E0B803011E82F6C6ABE861625 ) case (IDF2D2EFCFCAA060A180881D81395C002 ) I50BC02B32FFEA3FDDA09A1A76C72EDE6
: I72E47AC634CDDC2338CBBD5642F81090 = {16'h0000, I9C49DC380ED90CDC0B86D16428C58A39 }; I23CD01FB20FA1C856A43C90DA2FE8B37
: I72E47AC634CDDC2338CBBD5642F81090 = {16'h0003, IB733A674E6EDACC67D7A142D9C749704 , IE7811CA6D9DFDFCFDBDA2CB55876D5FC };
default : I72E47AC634CDDC2338CBBD5642F81090 = 32'b0; endcase else I72E47AC634CDDC2338CBBD5642F81090 = 32'b0; end
 always @(posedge ICCFB0F435B37370076102F325BC08D20 or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin if (~I9ED2A9117D3AEAF54CBA7AD69083BCB7 )
begin I9B8138DCE156F7C31EB5914EF01F183C <= 1'b0; IFFD0BAB32DEE73305A584A062E784936 <= 1'b1; I9C49DC380ED90CDC0B86D16428C58A39
<= {14'h0000, IDD2F1F37B45AD83BB6A8FD6BED814957 }; end else begin I9B8138DCE156F7C31EB5914EF01F183C <= (I9C49DC380ED90CDC0B86D16428C58A39 [1:0]
== 2'b00) ? 1'b1 : 1'b0; IFFD0BAB32DEE73305A584A062E784936 <= (I9C49DC380ED90CDC0B86D16428C58A39 [1:0] == 2'b11)
? 1'b1 : 1'b0; if (I7378609E0B803011E82F6C6ABE861625 & I684F27663FD8A3EFB4B2BC8B42792CD0 ) case (IDF2D2EFCFCAA060A180881D81395C002 )
I50BC02B32FFEA3FDDA09A1A76C72EDE6 : begin if (IE789C637CC57CC8ECB73F88C9790C5E4 [0]) I9C49DC380ED90CDC0B86D16428C58A39 [1:0]
<= I3C3096B9DAB1C65EA381C7E05B767FB3 [1:0]; end endcase end end endmodule 
 module IE63C8C66EC36AC972570F7B8665A4225 #( parameter I8F2F3EE9FE4B702742B51120C0EDA11A = 0, ID538F704AA7B227247264F05C613DABA
= 0, I394B9366718FFFBF01944193881668C1 = 0, I0A080290B2C86899F28748A119EE921C = 1 ) ( input wire ICCFB0F435B37370076102F325BC08D20 ,
input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire [11:0] I3D49ADB3C231E0C52B4EE7C42AB0DF8B , input wire
[3:0] IE789C637CC57CC8ECB73F88C9790C5E4 , input wire [31:0] I3C3096B9DAB1C65EA381C7E05B767FB3 , input wire I684F27663FD8A3EFB4B2BC8B42792CD0 ,
input wire I7378609E0B803011E82F6C6ABE861625 , input wire I6EC1BE4B18EC6AA3D88A5D45B614565E , output wire [2:0]
I42A419EB6EB8D11234AC3B2BCA0AE593 , output wire [2:0] IA41AC3CC6BC050DDC172724AB311315B , output wire [31:0] IB808853736ABE6034DB8E375F1F00E89
); `include "pcisig_constants.v"
 localparam [11:0] IB02BC4279E3AD90BA5C39FA16B9D5E8A = I8F2F3EE9FE4B702742B51120C0EDA11A ; localparam [11:0] IF594A0D212815344BE3693C306BF4EA2
= I8F2F3EE9FE4B702742B51120C0EDA11A + 12'h008; localparam [11:0] IDCC70C628E320A5251A1D0336068E6BB = I8F2F3EE9FE4B702742B51120C0EDA11A
+ 12'h00c; localparam [11:0] I87E36DB7D013BD93A24A5825D9370D13 = I8F2F3EE9FE4B702742B51120C0EDA11A + 12'h010; localparam
[3:0] I713C1A67C055ED94E63F28BD6B231361 = 4'h0; localparam [3:0] I81B2E848E59A16CC45F12458AC9C3755 = 4'b0001; localparam
[5:0] IBAB99C522164E1AC8426D8D04A5A59BA = 6'b000001; localparam [7:0] I3CFC8E9960B942C3792B7333D31D75D5 = ID538F704AA7B227247264F05C613DABA ;
localparam [3:0] I1D7F4405C57C37585B654ACB2055ED09 = I0A080290B2C86899F28748A119EE921C ;  reg [2:0] I2792804BC0B8F3DDCC1D08D4DE2F25DA ;
reg [2:0] IE763761FF58557F78DA03BEF9DCF712E ; reg [15:0] I009CBD7EE983A10185FB1BC848B106B8 ; reg [31:0] I72E47AC634CDDC2338CBBD5642F81090 ;
wire [11:0] IDF2D2EFCFCAA060A180881D81395C002 ;  assign I42A419EB6EB8D11234AC3B2BCA0AE593 = (I6EC1BE4B18EC6AA3D88A5D45B614565E )
? I2792804BC0B8F3DDCC1D08D4DE2F25DA : 3'b0; assign IA41AC3CC6BC050DDC172724AB311315B = (I6EC1BE4B18EC6AA3D88A5D45B614565E )
? IE763761FF58557F78DA03BEF9DCF712E : 3'b0; assign IB808853736ABE6034DB8E375F1F00E89 = I7378609E0B803011E82F6C6ABE861625
? I72E47AC634CDDC2338CBBD5642F81090 : 32'b0;  assign IDF2D2EFCFCAA060A180881D81395C002 = I3D49ADB3C231E0C52B4EE7C42AB0DF8B
& 12'hffc;  always @(*) begin if (I7378609E0B803011E82F6C6ABE861625 ) case (IDF2D2EFCFCAA060A180881D81395C002 )
IB02BC4279E3AD90BA5C39FA16B9D5E8A : I72E47AC634CDDC2338CBBD5642F81090 = {8'h0, I713C1A67C055ED94E63F28BD6B231361 ,
I1D7F4405C57C37585B654ACB2055ED09 , I3CFC8E9960B942C3792B7333D31D75D5 , IAD7735E1C92EEFA900A9BB537EC5BC75 }; IF594A0D212815344BE3693C306BF4EA2
: I72E47AC634CDDC2338CBBD5642F81090 = {16'b0, 1'b0, IE763761FF58557F78DA03BEF9DCF712E , 4'b0, I2792804BC0B8F3DDCC1D08D4DE2F25DA ,
5'b0}; IDCC70C628E320A5251A1D0336068E6BB :  I72E47AC634CDDC2338CBBD5642F81090 = (I394B9366718FFFBF01944193881668C1 )
? 32'h0003f012 : 32'h0003f011; I87E36DB7D013BD93A24A5825D9370D13 : I72E47AC634CDDC2338CBBD5642F81090 = 32'b0;  default :
I72E47AC634CDDC2338CBBD5642F81090 = 32'b0; endcase else I72E47AC634CDDC2338CBBD5642F81090 = 32'b0; end  always @(posedge
ICCFB0F435B37370076102F325BC08D20 or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin if (~I9ED2A9117D3AEAF54CBA7AD69083BCB7 )
begin I009CBD7EE983A10185FB1BC848B106B8 <= 16'b0; I2792804BC0B8F3DDCC1D08D4DE2F25DA <= 3'b0; IE763761FF58557F78DA03BEF9DCF712E
<= 3'b0; end else begin if (I7378609E0B803011E82F6C6ABE861625 & I684F27663FD8A3EFB4B2BC8B42792CD0 ) case (IDF2D2EFCFCAA060A180881D81395C002 )
IF594A0D212815344BE3693C306BF4EA2 : begin if (IE789C637CC57CC8ECB73F88C9790C5E4 [0]) I2792804BC0B8F3DDCC1D08D4DE2F25DA
<= I3C3096B9DAB1C65EA381C7E05B767FB3 [7:5]; if (IE789C637CC57CC8ECB73F88C9790C5E4 [1]) IE763761FF58557F78DA03BEF9DCF712E
<= I3C3096B9DAB1C65EA381C7E05B767FB3 [14:12]; end I87E36DB7D013BD93A24A5825D9370D13 : begin if (IE789C637CC57CC8ECB73F88C9790C5E4 [0])
begin I009CBD7EE983A10185FB1BC848B106B8 [1:0] <= I3C3096B9DAB1C65EA381C7E05B767FB3 [1:0];  I009CBD7EE983A10185FB1BC848B106B8 [3]
<= I3C3096B9DAB1C65EA381C7E05B767FB3 [3];  I009CBD7EE983A10185FB1BC848B106B8 [6] <= I3C3096B9DAB1C65EA381C7E05B767FB3 [6];
 end end endcase end end endmodule 
  module I2296FC491415818D18357D6C2D700C14 #( parameter IFC1FF746397E6A576E9FEB281890A248 = "NONE", IAF1DF965ED0D670C125D16FDF91B875B
= 0, IB7B379BA36F36F0638F4F33C7598CC85 = 0, ID9DCCEB6B5B42C479CB9D2B3C992035D = 1, I251C6E5612F7B344EC3156CB9A93BE5B
= "NONE", ID7A688D3DA9A2C539FE87FC8998248CB = 0, I96DBC3D130FB2B57DFB76E3E87DF89D2 = 1, I87B53E44EDBDCDA1796FB105323D3B17
= "NONE", IF9554E0938E353BDC05ABE0C628E3BE9 = 0, I37C708634F442A3B0568DA0BB576511F = 0, I7B125DA60401B7C86EB027E9E9262847
= 1, I8BEE88809FA5712893BC59FF0E17ADB2 = "NONE", I7DF5A90920A562D09AA22D2DFA657124 = 0, I0243B4A4E84E0712929C806F438E6AA9
= 1, I7050B96C0C45A812BBFC45C2A30F272C = "NONE", IB7C70D5D7B0DDF146F4D402BEE6F6FA6 = 0, I1CBD8B214B4765FBC7FA828F0C62BC94
= 0, I677BE3663880CBE6E5AE2C431F3FDD4D = 1, I1CF1EE9FA60C0CDB15DD404CC8A269E5 = "NONE", I34F020684BFF4B1EAA406E693751B71D
= 0, IFB94B817F0BC84EC0734110F6EDE475A = 1, I512A575E055CF9235066DBE4051242CB = 24'h000000, I391BF6A9C9F2ABEEA227F0E1F3F50A4F
= 16'h0000, IF0D7F78B99E50997A728E3731A197225 = 0, I9606837003EFA36A64A97C352D3D89A3 = "INTA", I4C1994114E1C49B9376320858F4E71F9
= 8'h00, I2CB8399B2A61CDA9DB269D3567018E65 = 16'h0000, I46C5269B9FB24EF04CE2CC341C288EC7 = 16'h0000, I3C9AD458B89B2FAABD743BF4E13BF421
= 16'h0000, I73ABD5619A9FB885445AC1E288EAF7F8 = 0, IBDE0431C8F903800F409661F4F56FD80 = 0, I394B9366718FFFBF01944193881668C1
= 0 ) ( input wire ICCFB0F435B37370076102F325BC08D20 , input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire
[31:0] ICB680FEAB46B6D635CD9DD6BB49A6A20 , input wire [31:0] I8FF768DAF4C56D1B2D217B2C02B6D4EC , input wire [31:0]
I9E5E6E86745F53F982BC3862031A206B , input wire [31:0] I3AD72E1D6C16169DB8A27F1681293009 , input wire [31:0] I0DE44F162EF92573C5DE1249527F6E9D ,
input wire [31:0] I2E9CC9AFC2E4742F852CB037CFC7E0A1 , input wire [63:0] I8B1798242C3B0E655181D0D365813614 , input
wire IE145222FDBDC80109E12FA72D3D3C655 , input wire ID43AC1009727D128F1C5DFE4640CA5AB , input wire IB610431939CB8180EAC2403672BAF58D ,
input wire [7:0] I3C7A9FA839F554D8898020C4831479E2 , input wire [4:0] I74A0936EE8FD1443A2C6745A4F3F6B5E , input
wire [2:0] I369BA2FFB5D41DF25F9BC3AB126D6607 , input wire [31:0] I1C0271AD5E8E9E9164909E468AD0B212 , input wire
I6EC1BE4B18EC6AA3D88A5D45B614565E , input wire I56148DDDF284443347FFCF4F9C3BE61A , input wire I24C403550AE065D7D1B7266142886226 ,
input wire [11:0] I438B8BD876741F9B46EB770E92F808B7 , input wire I5FE75BE614D4F52DB327549B36203350 , input wire
[31:0] I3D6C771D05CA1A769E61302C086494B8 , input wire [3:0] I357B3043EDACE3EBECE8F54D79B9F90A , input wire I0AAD559CF33A5CBA597990658774FEB3 ,
input wire I923204A95D8CBB206587CF32BEDCF4EF , output wire ICF9D8FD31DFC7D20DAF939C6D75F1518 , output wire IDF550B17734BF16B7E410B19BB31E276 ,
output wire I8ED9B9C1D9F58C5D06A9443AD901E8C6 , output wire IA976D63BEECA80DCE31365CF56EC0248 , output wire I5E3CE5AF5C34D232BFB139B63D9912B4 ,
output wire IBEF3E5F9395E2C7822AE03D6461DEBBB , output wire I7E6CFD6A7DCAB9CD2188D044C7D716A6 , output wire I3A34691662384260F0524DD7F650E75A ,
output wire IC2F58AB5028C1D2C53C6EF47A4975D0A , output wire [2:0] I112E0A79129A8BC6DD4C13647C31F8A0 , output wire
IE4B6DD43E04940631EF58BA04EA58997 , output wire I3A095084CDFDFA56A0E67616A78D3B25 , output wire I81CD7F184DF8D58A1F2324E975A6816C ,
output wire I83C4A4200EB2B3F6766D338284ECAAAF , output wire [2:0] I42A419EB6EB8D11234AC3B2BCA0AE593 , output wire
[2:0] IA41AC3CC6BC050DDC172724AB311315B , output wire I31CF69FF368B36B4D6612DF16B3ABC6B , output wire [31:0] IFE4A8CBA73734C6F0F0A078027E053D4 ,
output wire ID7A2A8B1E9D92B60194D5FAFAAB15208 , output wire IF274FAF97F5BACD693913BB418717A9D , output wire ID95C13E7EE1CFE6A8743FF9E62C25873 ,
output wire [10:0] IC58E411F24D810EF60A7B8638ABCC0BB , output wire I89CFFA73C7546481B72B0FB06D799AEE , output wire
I270ED686C2EF2C1C8B5B55EC4A5AAE84 , output wire ID5CCD4858CB5CC1B2EDEC682C7DE5AAD , output wire [31:0] I7D901091F9E0741061C75B54467D48A0
); `include "pcisig_constants.v"
 wire I528E34D2616570F6EB46E6E5A1689145 ; wire I5917F25EB5F020E0FEEB03EB956B3110 ; wire [11:0] IB49B50ED865F168D88C6EEBE96037C6E ;
wire [3:0] I183F148259060A23AC5E3DDBA1A409BD ; wire [31:0] I713670B3E894AB8B96764601F4FAD0A2 ; wire IBF48CFBD55119BD5D5AC0924CB673A2D ;
wire I8228086CD6BE873CD8E5EC62E459FEE8 ; wire IDAAB77FF78E6FA00D5A2E8600E96D156 ; wire I35A84B07F621AAD3B8596FBB41D3BB56 ;
wire I264580EA60DA3B2C5F03A620CFFC8AC8 ; wire IDAB3311066C56CFA851AD88D742521CC ; wire IA9369F8E522D76A4A2FB9CD46042A105 ;
wire IA1C5C4E78E2E56FD7177C302A7D223D4 ; wire I7ED71D3164ABC636AC5046B7E263FD03 ; wire [31:0] I6795B29551221467FFA6B7172DDA857D ;
wire IC0BDBEBC525B0F341D945F7586737805 ; wire I3048808F55068691CE04FEE2290AD354 ; wire I3A5FA9388628E5BE540E9EFA5A8A8AD0 ;
wire IF141F442E46E1CD59416531C214271F0 ; wire IB97F5BBF0732A355B8815AF36CD7C371 ; wire I39C3F8AA930CA6B1D9BC91786E27BC33 ;
wire I69BA038645155F12D6DFFF9C02EC3BE6 ; wire [31:0] ID9518A317572A0F59B950EF0E9602856 ; wire [5:0] IDDF260B92ADEBC1228A3C40D8F02ABB2 ;
wire [31:0] IBAD931958837224592F6A8D53ABD597B ; wire I88EAC02A1C9BA6648FAF51D1472253E6 ; wire IBA4050AD6F895B1AC3002D1A6C52B5FB ;
wire [31:0] I4FADCAEAE1DBE98C9FDAB11A1496AA63 ; wire [2:0] I6311EE8E4FBF32449E3D86CE286FFF12 ; wire [2:0] IDAF814B27DE872458FE905492366EC1F ;
wire [31:0] I3AFE1E2D1580EE3708616A828EEC91F9 ; wire [31:0] I4DF5B06333AF72835BFE083ACDE5B05B ; wire [31:0] I98308209671212A3C88A9644B503FA02 ;
wire IB4C822D6BFAE40F12254437B18142B8A ; wire I30157CAB406F288B630EF42C05ACC134 ; wire I82635882370B55739EA7454635CE3A41 ;
wire [10:0] IE38989B54E8F0643FD2DC5F4F7B5BCC6 ; wire I42E863B8B97EAE3620723BFD560E96F6 ; wire I5ADEE764CD8A8EACE17ED8F55EC633AC ;
wire I0E46034C0DD5EFC22C80F9C23EBDDCB7 ; wire [31:0] I7A347A14A6112DE258293F0AA5074560 ;  localparam [11:0] IA7EE8A611353335C5559FF1DB8FBF816
= (IF0D7F78B99E50997A728E3731A197225 ) ? I43C945338ADA718C47F9AC36AE9ADB8A : IC8E275CE62D6604F5CC30E6E067A1EA0 ;
 assign ICF9D8FD31DFC7D20DAF939C6D75F1518 = IC0BDBEBC525B0F341D945F7586737805 ; assign IDF550B17734BF16B7E410B19BB31E276
= I5917F25EB5F020E0FEEB03EB956B3110 ; assign I8ED9B9C1D9F58C5D06A9443AD901E8C6 = IDDF260B92ADEBC1228A3C40D8F02ABB2 [0];
assign IA976D63BEECA80DCE31365CF56EC0248 = IDDF260B92ADEBC1228A3C40D8F02ABB2 [1]; assign I5E3CE5AF5C34D232BFB139B63D9912B4
= IDDF260B92ADEBC1228A3C40D8F02ABB2 [2]; assign IBEF3E5F9395E2C7822AE03D6461DEBBB = IDDF260B92ADEBC1228A3C40D8F02ABB2 [3];
assign I7E6CFD6A7DCAB9CD2188D044C7D716A6 = IDDF260B92ADEBC1228A3C40D8F02ABB2 [4]; assign I3A34691662384260F0524DD7F650E75A
= IDDF260B92ADEBC1228A3C40D8F02ABB2 [5]; assign IC2F58AB5028C1D2C53C6EF47A4975D0A = (IDDF260B92ADEBC1228A3C40D8F02ABB2 )
? 1'b1 : 1'b0; assign I112E0A79129A8BC6DD4C13647C31F8A0 = (I528E34D2616570F6EB46E6E5A1689145 | IDDF260B92ADEBC1228A3C40D8F02ABB2 )
? I73ABD5619A9FB885445AC1E288EAF7F8 : 3'b0; assign IE4B6DD43E04940631EF58BA04EA58997 = I3048808F55068691CE04FEE2290AD354 ;
assign I3A095084CDFDFA56A0E67616A78D3B25 = I3A5FA9388628E5BE540E9EFA5A8A8AD0 ; assign I81CD7F184DF8D58A1F2324E975A6816C
= IF141F442E46E1CD59416531C214271F0 ; assign I83C4A4200EB2B3F6766D338284ECAAAF = IB97F5BBF0732A355B8815AF36CD7C371 ;
assign I42A419EB6EB8D11234AC3B2BCA0AE593 = I6311EE8E4FBF32449E3D86CE286FFF12 ; assign IA41AC3CC6BC050DDC172724AB311315B
= IDAF814B27DE872458FE905492366EC1F ; assign I31CF69FF368B36B4D6612DF16B3ABC6B = I88EAC02A1C9BA6648FAF51D1472253E6 ;
assign IFE4A8CBA73734C6F0F0A078027E053D4 = I98308209671212A3C88A9644B503FA02 ; assign ID7A2A8B1E9D92B60194D5FAFAAB15208
= IB4C822D6BFAE40F12254437B18142B8A ; assign IF274FAF97F5BACD693913BB418717A9D = I30157CAB406F288B630EF42C05ACC134 ;
assign ID95C13E7EE1CFE6A8743FF9E62C25873 = I82635882370B55739EA7454635CE3A41 ; assign IC58E411F24D810EF60A7B8638ABCC0BB
= IE38989B54E8F0643FD2DC5F4F7B5BCC6 ; assign I89CFFA73C7546481B72B0FB06D799AEE = I42E863B8B97EAE3620723BFD560E96F6 ;
assign I270ED686C2EF2C1C8B5B55EC4A5AAE84 = I5ADEE764CD8A8EACE17ED8F55EC633AC ; assign ID5CCD4858CB5CC1B2EDEC682C7DE5AAD
= I7ED71D3164ABC636AC5046B7E263FD03 ; assign I7D901091F9E0741061C75B54467D48A0 = I6795B29551221467FFA6B7172DDA857D ;
  assign I0E46034C0DD5EFC22C80F9C23EBDDCB7 = |I1C0271AD5E8E9E9164909E468AD0B212 ; assign I7A347A14A6112DE258293F0AA5074560
= ID9518A317572A0F59B950EF0E9602856 | IBAD931958837224592F6A8D53ABD597B | I4FADCAEAE1DBE98C9FDAB11A1496AA63 | I3AFE1E2D1580EE3708616A828EEC91F9
| I4DF5B06333AF72835BFE083ACDE5B05B ;  IC3C2C92E294852CA4AE110FD59776962 #( .IF0D7F78B99E50997A728E3731A197225 (IF0D7F78B99E50997A728E3731A197225 ),
.I73ABD5619A9FB885445AC1E288EAF7F8 (I73ABD5619A9FB885445AC1E288EAF7F8 ) ) IB420C4D1279F971E867FA537CA4D6E82 ( .ICCFB0F435B37370076102F325BC08D20
(ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .IE145222FDBDC80109E12FA72D3D3C655
(IE145222FDBDC80109E12FA72D3D3C655 ), .I369BA2FFB5D41DF25F9BC3AB126D6607 (I369BA2FFB5D41DF25F9BC3AB126D6607 ), .I8E073ABA74C317770ABA5D59E6FA0BFF
(IBA4050AD6F895B1AC3002D1A6C52B5FB ), .I3C3096B9DAB1C65EA381C7E05B767FB3 (I7A347A14A6112DE258293F0AA5074560 ), .I438B8BD876741F9B46EB770E92F808B7
(I438B8BD876741F9B46EB770E92F808B7 ), .I5FE75BE614D4F52DB327549B36203350 (I5FE75BE614D4F52DB327549B36203350 ), .I782B24592AE65A017A87162AE1B27668
(I3D6C771D05CA1A769E61302C086494B8 ), .I357B3043EDACE3EBECE8F54D79B9F90A (I357B3043EDACE3EBECE8F54D79B9F90A ), .I0AAD559CF33A5CBA597990658774FEB3
(I0AAD559CF33A5CBA597990658774FEB3 ), .I923204A95D8CBB206587CF32BEDCF4EF (I923204A95D8CBB206587CF32BEDCF4EF ), .I4A07557713C4283E634548A55A81AE55
(I528E34D2616570F6EB46E6E5A1689145 ), .IDF550B17734BF16B7E410B19BB31E276 (I5917F25EB5F020E0FEEB03EB956B3110 ), .I2E09014E801CDE025E646C14A7A88E8D
(IB49B50ED865F168D88C6EEBE96037C6E ), .I095F5745EA5D8A16BF789BA5B07338AA (I183F148259060A23AC5E3DDBA1A409BD ), .IB808853736ABE6034DB8E375F1F00E89
(I713670B3E894AB8B96764601F4FAD0A2 ), .I14BCC8E29270920B2D04C15BCF409C2F (IBF48CFBD55119BD5D5AC0924CB673A2D ), .I58DCF4F773FDA57377E940331963F6F2
(I8228086CD6BE873CD8E5EC62E459FEE8 ), .I34D5C55E6A7E8D35B8981814BB90440B (IDAAB77FF78E6FA00D5A2E8600E96D156 ), .ID7CE65853F1A17B2A146805CE598364F
(I35A84B07F621AAD3B8596FBB41D3BB56 ), .I207147984DF21E60B2451E00D7A06100 (I264580EA60DA3B2C5F03A620CFFC8AC8 ), .I25F92BF03720992A727F6B9F19ACA644
(IDAB3311066C56CFA851AD88D742521CC ), .I6A36AAB8630033974E1F982DFA8A6F7E (IA9369F8E522D76A4A2FB9CD46042A105 ), .I8B94BE4224AE909FF34FA01D95C810CE
(IA1C5C4E78E2E56FD7177C302A7D223D4 ), .ID5CCD4858CB5CC1B2EDEC682C7DE5AAD (I7ED71D3164ABC636AC5046B7E263FD03 ), .I6E43903839286F6F3DAB2A247E5C3D77
(I6795B29551221467FFA6B7172DDA857D ) ); ID6D6E4DEEE2F225D2FE2E68AEDBFADC7 #( .I9449A4DEE4C71770D9A5095574AED415
(I8125345218ED2F68A2205656CAD621A2 ), .I4700AD5A2ED246219F585C312B2124C9 (I512A575E055CF9235066DBE4051242CB ), .IB2FE05230F3A440BAF4BE98DCA56829F
(I391BF6A9C9F2ABEEA227F0E1F3F50A4F ), .I28B2C4B454208AC784C97EA8274B9503 (IF0D7F78B99E50997A728E3731A197225 ), .I7F482C6D7FFF305AD90ABABC0457155E
(I9606837003EFA36A64A97C352D3D89A3 ), .IBDE0431C8F903800F409661F4F56FD80 (IBDE0431C8F903800F409661F4F56FD80 ), .IE0E04F5EA496E6FD62B9A6B66E33F418
(I4C1994114E1C49B9376320858F4E71F9 ), .I060C01BCB8E6DC3D4B74BEFA66D56545 (I2CB8399B2A61CDA9DB269D3567018E65 ), .ID34BC6EE8891CF37121D63EE0EAD6385
(I46C5269B9FB24EF04CE2CC341C288EC7 ), .I9831646508922ACBA52B47759E0BAD32 (I3C9AD458B89B2FAABD743BF4E13BF421 ) )
I617CBE084F8475F4DC0DA892B8855F84 ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .I1C0271AD5E8E9E9164909E468AD0B212 (I0E46034C0DD5EFC22C80F9C23EBDDCB7 ), .I9119CE851F731CBC5834D0370CCA6908
(I88EAC02A1C9BA6648FAF51D1472253E6 ), .I3D49ADB3C231E0C52B4EE7C42AB0DF8B (IB49B50ED865F168D88C6EEBE96037C6E ), .IE789C637CC57CC8ECB73F88C9790C5E4
(I183F148259060A23AC5E3DDBA1A409BD ), .I3C3096B9DAB1C65EA381C7E05B767FB3 (I713670B3E894AB8B96764601F4FAD0A2 ), .I684F27663FD8A3EFB4B2BC8B42792CD0
(IBF48CFBD55119BD5D5AC0924CB673A2D ), .I7378609E0B803011E82F6C6ABE861625 (IA1C5C4E78E2E56FD7177C302A7D223D4 ), .ICF9D8FD31DFC7D20DAF939C6D75F1518
(IC0BDBEBC525B0F341D945F7586737805 ), .IE4B6DD43E04940631EF58BA04EA58997 (I3048808F55068691CE04FEE2290AD354 ), .I3A095084CDFDFA56A0E67616A78D3B25
(I3A5FA9388628E5BE540E9EFA5A8A8AD0 ), .I81CD7F184DF8D58A1F2324E975A6816C (IF141F442E46E1CD59416531C214271F0 ), .I83C4A4200EB2B3F6766D338284ECAAAF
(IB97F5BBF0732A355B8815AF36CD7C371 ), .IDA2B8A1BA5BD091F8C569BAA1CE5FED0 (I39C3F8AA930CA6B1D9BC91786E27BC33 ), .I9AFDACCEB4D156D714A2B8E72990FDA6
(I69BA038645155F12D6DFFF9C02EC3BE6 ), .IB808853736ABE6034DB8E375F1F00E89 (ID9518A317572A0F59B950EF0E9602856 ) );
I7649039BBE19689793FEE4FADDDEF1E8 #( .IFDFBBCC4A729BEC2BC4A96ABA6A686B0 (IAF1DF965ED0D670C125D16FDF91B875B ), .I60C4892BECCA6E2B2FE143BD923A22CA
(IF9554E0938E353BDC05ABE0C628E3BE9 ), .I614E1E615DEE042F64BC57A314245927 (IB7C70D5D7B0DDF146F4D402BEE6F6FA6 ), .I2E554B9CAB59E598058B7921DA36D560
(IFC1FF746397E6A576E9FEB281890A248 ), .I259BF2DBCEAAB39C062C08519379767E (IB7B379BA36F36F0638F4F33C7598CC85 ), .I2B0035459578DEB60AE2E24DF687E762
(ID9DCCEB6B5B42C479CB9D2B3C992035D ), .IB04EEBB96EE0ED06EDBB60ACE60A4A93 (I251C6E5612F7B344EC3156CB9A93BE5B ), .I86027F65FEA0494C8A49DAFE67EDAE13
(ID7A688D3DA9A2C539FE87FC8998248CB ), .ID3FF77989ABAC7B0FC1DE518FA7D21E6 (I96DBC3D130FB2B57DFB76E3E87DF89D2 ), .IDD5BBB6DF3D487FCF2DA81CA8794849C
(I87B53E44EDBDCDA1796FB105323D3B17 ), .I4E3CEE40D32239479A1163B2D85B5FA7 (I37C708634F442A3B0568DA0BB576511F ), .I41D8D6036479734032C1711509A67D83
(I7B125DA60401B7C86EB027E9E9262847 ), .I0AA7FFBF9C00DEF85FA40AFFAF675794 (I8BEE88809FA5712893BC59FF0E17ADB2 ), .I6104B7636177E429318BE1C790C3CB49
(I7DF5A90920A562D09AA22D2DFA657124 ), .I0D8F74FCCB77AD67CAB98890C8885156 (I0243B4A4E84E0712929C806F438E6AA9 ), .IFB616CA07D005C26A9BA5823D543CCBD
(I7050B96C0C45A812BBFC45C2A30F272C ), .IA67F3F71E4F9434D68536978B81F91DA (I1CBD8B214B4765FBC7FA828F0C62BC94 ), .IB6ECC5AF80982DE8999481CA0E9A481A
(I677BE3663880CBE6E5AE2C431F3FDD4D ), .I21FC0FBCD63A328488B305A90691197D (I1CF1EE9FA60C0CDB15DD404CC8A269E5 ), .I02E3D3076327F179BFEC2E663B0EAE70
(I34F020684BFF4B1EAA406E693751B71D ), .I6D6B05AA28D91BF74A2607970B27F65D (IFB94B817F0BC84EC0734110F6EDE475A ) )
I1A907F2B09600B273EEF91F54930FBC2 ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .I7195780B6CCA660A6833F98360035D81 (I8B1798242C3B0E655181D0D365813614 [63:32]),
.I077B3A3A6F38E8073B18F35643BD4B02 (I8B1798242C3B0E655181D0D365813614 [31:0]), .I660A2BFC1099D715D966FB7D0E899778
(I8228086CD6BE873CD8E5EC62E459FEE8 ), .I52BCA73A227659ABF278B7B041C2D33A (IDAAB77FF78E6FA00D5A2E8600E96D156 ), .I275F5F6495E251A9F1E0A46729B18393
(I35A84B07F621AAD3B8596FBB41D3BB56 ), .ICB680FEAB46B6D635CD9DD6BB49A6A20 (ICB680FEAB46B6D635CD9DD6BB49A6A20 ), .I8FF768DAF4C56D1B2D217B2C02B6D4EC
(I8FF768DAF4C56D1B2D217B2C02B6D4EC ), .I9E5E6E86745F53F982BC3862031A206B (I9E5E6E86745F53F982BC3862031A206B ), .I3AD72E1D6C16169DB8A27F1681293009
(I3AD72E1D6C16169DB8A27F1681293009 ), .I0DE44F162EF92573C5DE1249527F6E9D (I0DE44F162EF92573C5DE1249527F6E9D ), .I2E9CC9AFC2E4742F852CB037CFC7E0A1
(I2E9CC9AFC2E4742F852CB037CFC7E0A1 ), .I003A2455D9D9F27B56BE4B6A6E330845 (I39C3F8AA930CA6B1D9BC91786E27BC33 ), .I61583F0AD8ACE3D2B571B36EFC23311D
(I69BA038645155F12D6DFFF9C02EC3BE6 ), .I332C3203B01AAFA54A288D09DDEB7AFB (ID43AC1009727D128F1C5DFE4640CA5AB ), .I3D2849BFA4C1331FDDB8A39BF571CD91
(IB610431939CB8180EAC2403672BAF58D ), .I6E16E1B891ED18DC65EFF37952418F3C (IB49B50ED865F168D88C6EEBE96037C6E [2]),
.I410A0939BF5AB6CE2A725DB6210E101F (I713670B3E894AB8B96764601F4FAD0A2 ), .I22B24791BA0E7AA2C686B1B2D776C636 (IBF48CFBD55119BD5D5AC0924CB673A2D ),
.IAF378590D5A80382A321B73D17E05142 (IDDF260B92ADEBC1228A3C40D8F02ABB2 ), .IDCFC89CB36B3EFB6258338EC62FFDD79 (IBAD931958837224592F6A8D53ABD597B )
); IF44E5E7AB65AFFA1AF3DA949DB91C839 #( .I8F2F3EE9FE4B702742B51120C0EDA11A (I8125345218ED2F68A2205656CAD621A2 ),
.ID538F704AA7B227247264F05C613DABA (IA7EE8A611353335C5559FF1DB8FBF816 ) ) I191AE9CE91C1B22E4AE2BF8631B30918 ( .ICCFB0F435B37370076102F325BC08D20
(ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .I3D49ADB3C231E0C52B4EE7C42AB0DF8B
(IB49B50ED865F168D88C6EEBE96037C6E ), .IE789C637CC57CC8ECB73F88C9790C5E4 (I183F148259060A23AC5E3DDBA1A409BD ), .I3C3096B9DAB1C65EA381C7E05B767FB3
(I713670B3E894AB8B96764601F4FAD0A2 ), .I684F27663FD8A3EFB4B2BC8B42792CD0 (IBF48CFBD55119BD5D5AC0924CB673A2D ), .I7378609E0B803011E82F6C6ABE861625
(IA9369F8E522D76A4A2FB9CD46042A105 ), .I31CF69FF368B36B4D6612DF16B3ABC6B (I88EAC02A1C9BA6648FAF51D1472253E6 ), .I26F316E89E4B007444B724CD95758235
(IBA4050AD6F895B1AC3002D1A6C52B5FB ), .IB808853736ABE6034DB8E375F1F00E89 (I4FADCAEAE1DBE98C9FDAB11A1496AA63 ) );
IE63C8C66EC36AC972570F7B8665A4225 #( .I8F2F3EE9FE4B702742B51120C0EDA11A (IC8E275CE62D6604F5CC30E6E067A1EA0 ), .ID538F704AA7B227247264F05C613DABA
(0), .I394B9366718FFFBF01944193881668C1 (I394B9366718FFFBF01944193881668C1 ), .I0A080290B2C86899F28748A119EE921C
(1) ) I2A3F2A5CBC5AE0DD0620353468BA1D81 ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ),
.I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .I3D49ADB3C231E0C52B4EE7C42AB0DF8B (IB49B50ED865F168D88C6EEBE96037C6E ),
.IE789C637CC57CC8ECB73F88C9790C5E4 (I183F148259060A23AC5E3DDBA1A409BD ), .I3C3096B9DAB1C65EA381C7E05B767FB3 (I713670B3E894AB8B96764601F4FAD0A2 ),
.I684F27663FD8A3EFB4B2BC8B42792CD0 (IBF48CFBD55119BD5D5AC0924CB673A2D ), .I7378609E0B803011E82F6C6ABE861625 (IDAB3311066C56CFA851AD88D742521CC ),
.I6EC1BE4B18EC6AA3D88A5D45B614565E (I6EC1BE4B18EC6AA3D88A5D45B614565E ), .I42A419EB6EB8D11234AC3B2BCA0AE593 (I6311EE8E4FBF32449E3D86CE286FFF12 ),
.IA41AC3CC6BC050DDC172724AB311315B (IDAF814B27DE872458FE905492366EC1F ), .IB808853736ABE6034DB8E375F1F00E89 (I3AFE1E2D1580EE3708616A828EEC91F9 )
); generate if (IF0D7F78B99E50997A728E3731A197225 ) IB692DAE41499E4B01D446B8B28C804EB #( .I8F2F3EE9FE4B702742B51120C0EDA11A
(I43C945338ADA718C47F9AC36AE9ADB8A ), .I73ABD5619A9FB885445AC1E288EAF7F8 (I73ABD5619A9FB885445AC1E288EAF7F8 ), .I28B2C4B454208AC784C97EA8274B9503
(IF0D7F78B99E50997A728E3731A197225 ), .ID538F704AA7B227247264F05C613DABA (IC8E275CE62D6604F5CC30E6E067A1EA0 ) )
I39D757619EF5DEA91CD3A2B7CE5AFB30 ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .I3C7A9FA839F554D8898020C4831479E2 (I3C7A9FA839F554D8898020C4831479E2 ), .I74A0936EE8FD1443A2C6745A4F3F6B5E
(I74A0936EE8FD1443A2C6745A4F3F6B5E ), .I1C0271AD5E8E9E9164909E468AD0B212 (I1C0271AD5E8E9E9164909E468AD0B212 ), .I3D49ADB3C231E0C52B4EE7C42AB0DF8B
(IB49B50ED865F168D88C6EEBE96037C6E ), .IE789C637CC57CC8ECB73F88C9790C5E4 (I183F148259060A23AC5E3DDBA1A409BD ), .I3C3096B9DAB1C65EA381C7E05B767FB3
(I713670B3E894AB8B96764601F4FAD0A2 ), .I684F27663FD8A3EFB4B2BC8B42792CD0 (IBF48CFBD55119BD5D5AC0924CB673A2D ), .I7378609E0B803011E82F6C6ABE861625
(I264580EA60DA3B2C5F03A620CFFC8AC8 ), .I56148DDDF284443347FFCF4F9C3BE61A (I56148DDDF284443347FFCF4F9C3BE61A ), .I24C403550AE065D7D1B7266142886226
(I24C403550AE065D7D1B7266142886226 ), .IB808853736ABE6034DB8E375F1F00E89 (I4DF5B06333AF72835BFE083ACDE5B05B ), .IFE4A8CBA73734C6F0F0A078027E053D4
(I98308209671212A3C88A9644B503FA02 ), .ID7A2A8B1E9D92B60194D5FAFAAB15208 (IB4C822D6BFAE40F12254437B18142B8A ), .IF274FAF97F5BACD693913BB418717A9D
(I30157CAB406F288B630EF42C05ACC134 ), .ID95C13E7EE1CFE6A8743FF9E62C25873 (I82635882370B55739EA7454635CE3A41 ), .IC58E411F24D810EF60A7B8638ABCC0BB
(IE38989B54E8F0643FD2DC5F4F7B5BCC6 ), .I89CFFA73C7546481B72B0FB06D799AEE (I42E863B8B97EAE3620723BFD560E96F6 ), .I270ED686C2EF2C1C8B5B55EC4A5AAE84
(I5ADEE764CD8A8EACE17ED8F55EC633AC ) ); else begin assign I4DF5B06333AF72835BFE083ACDE5B05B = 32'b0; assign I98308209671212A3C88A9644B503FA02
= 32'b0; assign IB4C822D6BFAE40F12254437B18142B8A = 1'b0; assign I30157CAB406F288B630EF42C05ACC134 = 1'b0; assign
I82635882370B55739EA7454635CE3A41 = 1'b0; assign IE38989B54E8F0643FD2DC5F4F7B5BCC6 = 11'b0; assign I42E863B8B97EAE3620723BFD560E96F6
= 1'b0; assign I5ADEE764CD8A8EACE17ED8F55EC633AC = 1'b0; end endgenerate endmodule 
  module IF8888DF840520FCED3157D151D128B3B #( parameter IE50492CEE03959C13AD5E521CC7F2FEF = 0, I0B3C14F69FAC563649E26679A3D8B1CD
= 0, IFA272F301A5935EE15CB134524665363 = 0, IE690B7723F136DA02896C0728DDADB49 = 0, I55BE27080C370AF723A4FE096014E875
= 0, IB2560D175E4507798B84D6E659FD6373 = 0, I25B649490B20A1FEC9A1AA60AB0C6D5E = 0 ) ( input wire ICCFB0F435B37370076102F325BC08D20 ,
input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire IE145222FDBDC80109E12FA72D3D3C655 , input wire I2AD6292CA4A68298ECB0EB04E60DC338 ,
input wire I7E1B3386EACDCC0730096B4BEBD3FC11 , input wire IE10AAAB7732A262D17819D08F8A724BC , input wire IDF7BAD8C79D202960378A7387FEE4794 ,
input wire I57990336F36AA63E9FBA5533A4E25FA3 , input wire IED35F37F7AD8CD8C1B242C9C79E11FA3 , input wire [7:0] ID2BF5B6DEE97B309004C8AC7C3F5B8B3 ,
input wire [7:0] I3C7A9FA839F554D8898020C4831479E2 , input wire [4:0] I74A0936EE8FD1443A2C6745A4F3F6B5E , input
wire [2:0] I369BA2FFB5D41DF25F9BC3AB126D6607 , input wire [7:0] I2CB69D0EFAF8ADA6B6211F64BA9D2B52 , input wire [7:0]
I3EEF1AC61F6E4A2B704EBA11EF949965 , input wire [7:0] I25EC384599199AF35E4D0B3B873187EF , input wire [7:0] I8F57B8D98905C89F4D3B91CA626C25BA ,
input wire I56148DDDF284443347FFCF4F9C3BE61A , input wire I24C403550AE065D7D1B7266142886226 , input wire I5FE75BE614D4F52DB327549B36203350 ,
input wire I0AAD559CF33A5CBA597990658774FEB3 , input wire I923204A95D8CBB206587CF32BEDCF4EF , output wire I20CD33DEFBDF51E2A5352736B083738D ,
output wire I8ED9B9C1D9F58C5D06A9443AD901E8C6 , output wire IA976D63BEECA80DCE31365CF56EC0248 , output wire I5E3CE5AF5C34D232BFB139B63D9912B4 ,
output wire IBEF3E5F9395E2C7822AE03D6461DEBBB , output wire I7E6CFD6A7DCAB9CD2188D044C7D716A6 , output wire I3A34691662384260F0524DD7F650E75A ,
output wire [7:0] IC2F58AB5028C1D2C53C6EF47A4975D0A , output wire [7:0] ID3E7F4B58943229FEE6313A36B3F8693 , output
wire [4:0] I1FDEC1735547330C00A0B8DFE1FB10C3 , output wire I439AF6D496491F5F7C23217209B43C31 , output wire [31:0]
IFE4A8CBA73734C6F0F0A078027E053D4 , output wire ID7A2A8B1E9D92B60194D5FAFAAB15208 , output wire IF274FAF97F5BACD693913BB418717A9D ,
output wire ID95C13E7EE1CFE6A8743FF9E62C25873 , output wire I0DA874BD2204FA5231F61AC696D6584A , output wire I270ED686C2EF2C1C8B5B55EC4A5AAE84
); `include "pcisig_constants.v"
 localparam IBE3FC19439FEC0073D66B4DAC2FECC32 = 4'b0000, I310264643E51C96BF8FECF37C2EB7553 = 4'b0001, IAFB2BC0EA796EA2F143B022C32D56FCC
= 4'b0010, IB096F3B4C49EC3A522650D9969041D46 = 4'b0011, IA7E2C061B23F9C2D79751962637FF9F8 = 4'b0100, I02DAFFFA7BA0DF9723298CABE1A6EDF3
= 4'b0101, I0FBF38AB1DE3B938794F64EFEB6EEF04 = 4'b0110, I2512657214BD8CD9D7C9E46341FB6960 = 4'b0111, IA4F9276F2E3EF93B14F2B0FF3B2DDE74
= 4'b1000, I3AEAA310DC2EB1E6D2E2AB4DD0417BA2 = 4'b1001, I9CFCF3FC76F8BCD4AA7E722E67E01A89 = 4'b1010, IDA65D1282C0B7B2A86436F0450F882A3
= 4'b1011, I17BD3A950F8A3CC40AA8CA373AA26A5C = 4'b1100;  reg IDC8BCCAF6838A741E22C5D6213BD93DB ; reg IBB1C5765B30D0AAF14E2AF3F0F61A696 ;
reg I7CFDA4B8CD4F017B34A458F2130F1F2C ; reg I040F45C8B8CD2190DF8565751E1452CA ; reg IA0CE7A5E72A820959466307C122813D9 ;
reg IC2D075CC3D156038468427C3B77FAFCE ; reg I60C05F870B32C61B7CE3F165C499FB12 ; reg [7:0] I26AD306F3EB5A0DD0DA30F04952A3EF8 ;
reg [7:0] I7E9516402D6933186513EB5B37336278 ; reg [4:0] IA1EA4D4C05E159614ABC1E6D9CABE3BB ; reg [3:0] I91047088394D6A4116575942899FC337 ;
reg [3:0] ICBC89A2A67F0564ABA5BC46C474021BD ; reg [7:0] I6B25926923BB34891F18EDE430675796 ; reg [3:0] ID2E840891AA711130477F703743EDCF7 ;
reg I6D75F828BC25A6E4A9A4E45BE2A20DA5 ; reg ID038E78CE0FF71E71ACCE3E261678383 ; reg I9D1C45A4D6256BE0229612FD8C39AFBA ;
reg I31761EA46D336BB6B89BCC04E58CA62D ; reg IB97EB95EF3D656CF774FCC82AC2AE0FF ; reg [31:0] ID0A5ECECBEC8CE692F380DDF069E842F ;
reg I1877CB8174894BB7A9732E91A1794AAA ; reg [3:0] I7E04E8229BE60B48AAE3E1EB6511163A ; reg [3:0] ID22BB0550BCC1515614C8142FADDA171 ;
reg I612E93B17FEB6E7AE6FD9448B52CA816 ; reg I8D181359467F27637239CDAEE8A2F45A ;  assign I20CD33DEFBDF51E2A5352736B083738D
= IDC8BCCAF6838A741E22C5D6213BD93DB ; assign I8ED9B9C1D9F58C5D06A9443AD901E8C6 = IBB1C5765B30D0AAF14E2AF3F0F61A696 ;
assign IA976D63BEECA80DCE31365CF56EC0248 = I7CFDA4B8CD4F017B34A458F2130F1F2C ; assign I5E3CE5AF5C34D232BFB139B63D9912B4
= I040F45C8B8CD2190DF8565751E1452CA ; assign IBEF3E5F9395E2C7822AE03D6461DEBBB = IA0CE7A5E72A820959466307C122813D9 ;
assign I7E6CFD6A7DCAB9CD2188D044C7D716A6 = IC2D075CC3D156038468427C3B77FAFCE ; assign I3A34691662384260F0524DD7F650E75A
= I60C05F870B32C61B7CE3F165C499FB12 ; assign IC2F58AB5028C1D2C53C6EF47A4975D0A = I26AD306F3EB5A0DD0DA30F04952A3EF8 ;
assign ID3E7F4B58943229FEE6313A36B3F8693 = I7E9516402D6933186513EB5B37336278 ; assign I1FDEC1735547330C00A0B8DFE1FB10C3
= IA1EA4D4C05E159614ABC1E6D9CABE3BB ; assign I439AF6D496491F5F7C23217209B43C31 = IB97EB95EF3D656CF774FCC82AC2AE0FF ;
assign IFE4A8CBA73734C6F0F0A078027E053D4 = ID0A5ECECBEC8CE692F380DDF069E842F ; assign ID7A2A8B1E9D92B60194D5FAFAAB15208
= I1877CB8174894BB7A9732E91A1794AAA ; assign IF274FAF97F5BACD693913BB418717A9D = I612E93B17FEB6E7AE6FD9448B52CA816 ;
assign ID95C13E7EE1CFE6A8743FF9E62C25873 = (I7E04E8229BE60B48AAE3E1EB6511163A == I310264643E51C96BF8FECF37C2EB7553 )
? 1'b1 : 1'b0; assign I0DA874BD2204FA5231F61AC696D6584A = (I7E04E8229BE60B48AAE3E1EB6511163A == I17BD3A950F8A3CC40AA8CA373AA26A5C )
? 1'b1 : 1'b0; assign I270ED686C2EF2C1C8B5B55EC4A5AAE84 = I8D181359467F27637239CDAEE8A2F45A ;  always @(I91047088394D6A4116575942899FC337
or I7E04E8229BE60B48AAE3E1EB6511163A or I56148DDDF284443347FFCF4F9C3BE61A or I24C403550AE065D7D1B7266142886226 )
begin ID22BB0550BCC1515614C8142FADDA171 = I7E04E8229BE60B48AAE3E1EB6511163A ; case (I7E04E8229BE60B48AAE3E1EB6511163A )
IBE3FC19439FEC0073D66B4DAC2FECC32 : begin if ((|I91047088394D6A4116575942899FC337 ) & ~I56148DDDF284443347FFCF4F9C3BE61A )
ID22BB0550BCC1515614C8142FADDA171 = I310264643E51C96BF8FECF37C2EB7553 ; end I310264643E51C96BF8FECF37C2EB7553 :
begin if (I56148DDDF284443347FFCF4F9C3BE61A ) ID22BB0550BCC1515614C8142FADDA171 = IAFB2BC0EA796EA2F143B022C32D56FCC ;
end IAFB2BC0EA796EA2F143B022C32D56FCC : begin ID22BB0550BCC1515614C8142FADDA171 = IB096F3B4C49EC3A522650D9969041D46 ;
end IB096F3B4C49EC3A522650D9969041D46 : begin if (I6B25926923BB34891F18EDE430675796 == I9E0B4C1FB5C57E21C6F98D25B6A3CC40 )
ID22BB0550BCC1515614C8142FADDA171 = I17BD3A950F8A3CC40AA8CA373AA26A5C ; else ID22BB0550BCC1515614C8142FADDA171 =
IA7E2C061B23F9C2D79751962637FF9F8 ; end IA7E2C061B23F9C2D79751962637FF9F8 : begin ID22BB0550BCC1515614C8142FADDA171
= I0FBF38AB1DE3B938794F64EFEB6EEF04 ; end I0FBF38AB1DE3B938794F64EFEB6EEF04 : begin ID22BB0550BCC1515614C8142FADDA171
= I2512657214BD8CD9D7C9E46341FB6960 ; end I2512657214BD8CD9D7C9E46341FB6960 : begin ID22BB0550BCC1515614C8142FADDA171
= IA4F9276F2E3EF93B14F2B0FF3B2DDE74 ; end IA4F9276F2E3EF93B14F2B0FF3B2DDE74 : begin ID22BB0550BCC1515614C8142FADDA171
= I3AEAA310DC2EB1E6D2E2AB4DD0417BA2 ; end I3AEAA310DC2EB1E6D2E2AB4DD0417BA2 : begin ID22BB0550BCC1515614C8142FADDA171
= I9CFCF3FC76F8BCD4AA7E722E67E01A89 ; end I9CFCF3FC76F8BCD4AA7E722E67E01A89 : begin ID22BB0550BCC1515614C8142FADDA171
= IDA65D1282C0B7B2A86436F0450F882A3 ; end IDA65D1282C0B7B2A86436F0450F882A3 : begin if (I24C403550AE065D7D1B7266142886226 )
ID22BB0550BCC1515614C8142FADDA171 = IBE3FC19439FEC0073D66B4DAC2FECC32 ; end I17BD3A950F8A3CC40AA8CA373AA26A5C :
begin ID22BB0550BCC1515614C8142FADDA171 = IBE3FC19439FEC0073D66B4DAC2FECC32 ; end default : begin end endcase end
 always @(posedge ICCFB0F435B37370076102F325BC08D20 or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin if (~I9ED2A9117D3AEAF54CBA7AD69083BCB7 )
begin IDC8BCCAF6838A741E22C5D6213BD93DB <= 1'b0; IBB1C5765B30D0AAF14E2AF3F0F61A696 <= 1'b0; I7CFDA4B8CD4F017B34A458F2130F1F2C
<= 1'b0; I040F45C8B8CD2190DF8565751E1452CA <= 1'b0; IA0CE7A5E72A820959466307C122813D9 <= 1'b0; IC2D075CC3D156038468427C3B77FAFCE
<= 1'b0; I60C05F870B32C61B7CE3F165C499FB12 <= 1'b0; I26AD306F3EB5A0DD0DA30F04952A3EF8 <= 8'b0; I7E9516402D6933186513EB5B37336278
<= 8'b0; IA1EA4D4C05E159614ABC1E6D9CABE3BB <= 5'b0; I91047088394D6A4116575942899FC337 <= 4'b0; I6B25926923BB34891F18EDE430675796
<= 8'b0; ID2E840891AA711130477F703743EDCF7 <= 4'b0; ICBC89A2A67F0564ABA5BC46C474021BD <= 4'b0; I6D75F828BC25A6E4A9A4E45BE2A20DA5
<= 1'b0; ID038E78CE0FF71E71ACCE3E261678383 <= 1'b0; I9D1C45A4D6256BE0229612FD8C39AFBA <= 1'b0; I31761EA46D336BB6B89BCC04E58CA62D
<= 1'b0; IB97EB95EF3D656CF774FCC82AC2AE0FF <= 1'b0; ID0A5ECECBEC8CE692F380DDF069E842F <= 32'b0; I1877CB8174894BB7A9732E91A1794AAA
<= 1'b0; I7E04E8229BE60B48AAE3E1EB6511163A <= IBE3FC19439FEC0073D66B4DAC2FECC32 ; I612E93B17FEB6E7AE6FD9448B52CA816
<= 1'b0; I8D181359467F27637239CDAEE8A2F45A <= 1'b0; end else begin IB97EB95EF3D656CF774FCC82AC2AE0FF <= 1'b1; IDC8BCCAF6838A741E22C5D6213BD93DB
<= ((I369BA2FFB5D41DF25F9BC3AB126D6607 == 3'b000) ? IE145222FDBDC80109E12FA72D3D3C655 : 1'b0) | (((I369BA2FFB5D41DF25F9BC3AB126D6607
== 3'b001) && IE50492CEE03959C13AD5E521CC7F2FEF ) ? IE145222FDBDC80109E12FA72D3D3C655 : 1'b0) | (((I369BA2FFB5D41DF25F9BC3AB126D6607
== 3'b010) && I0B3C14F69FAC563649E26679A3D8B1CD ) ? IE145222FDBDC80109E12FA72D3D3C655 : 1'b0) | (((I369BA2FFB5D41DF25F9BC3AB126D6607
== 3'b011) && IFA272F301A5935EE15CB134524665363 ) ? IE145222FDBDC80109E12FA72D3D3C655 : 1'b0) | (((I369BA2FFB5D41DF25F9BC3AB126D6607
== 3'b100) && IE690B7723F136DA02896C0728DDADB49 ) ? IE145222FDBDC80109E12FA72D3D3C655 : 1'b0) | (((I369BA2FFB5D41DF25F9BC3AB126D6607
== 3'b101) && I55BE27080C370AF723A4FE096014E875 ) ? IE145222FDBDC80109E12FA72D3D3C655 : 1'b0) | (((I369BA2FFB5D41DF25F9BC3AB126D6607
== 3'b110) && IB2560D175E4507798B84D6E659FD6373 ) ? IE145222FDBDC80109E12FA72D3D3C655 : 1'b0) | (((I369BA2FFB5D41DF25F9BC3AB126D6607
== 3'b111) && I25B649490B20A1FEC9A1AA60AB0C6D5E ) ? IE145222FDBDC80109E12FA72D3D3C655 : 1'b0); IBB1C5765B30D0AAF14E2AF3F0F61A696
<= I2AD6292CA4A68298ECB0EB04E60DC338 ; I7CFDA4B8CD4F017B34A458F2130F1F2C <= I7E1B3386EACDCC0730096B4BEBD3FC11 ;
I040F45C8B8CD2190DF8565751E1452CA <= IE10AAAB7732A262D17819D08F8A724BC ; IA0CE7A5E72A820959466307C122813D9 <= IDF7BAD8C79D202960378A7387FEE4794 ;
IC2D075CC3D156038468427C3B77FAFCE <= I57990336F36AA63E9FBA5533A4E25FA3 ; I60C05F870B32C61B7CE3F165C499FB12 <= IED35F37F7AD8CD8C1B242C9C79E11FA3 ;
I26AD306F3EB5A0DD0DA30F04952A3EF8 <= ID2BF5B6DEE97B309004C8AC7C3F5B8B3 ; I91047088394D6A4116575942899FC337 <= ID2E840891AA711130477F703743EDCF7
^ ICBC89A2A67F0564ABA5BC46C474021BD ; ID2E840891AA711130477F703743EDCF7 <= {I31761EA46D336BB6B89BCC04E58CA62D ,
I9D1C45A4D6256BE0229612FD8C39AFBA , ID038E78CE0FF71E71ACCE3E261678383 , I6D75F828BC25A6E4A9A4E45BE2A20DA5 }; I6D75F828BC25A6E4A9A4E45BE2A20DA5
<= |I2CB69D0EFAF8ADA6B6211F64BA9D2B52 ; ID038E78CE0FF71E71ACCE3E261678383 <= |I3EEF1AC61F6E4A2B704EBA11EF949965 ;
I9D1C45A4D6256BE0229612FD8C39AFBA <= |I25EC384599199AF35E4D0B3B873187EF ; I31761EA46D336BB6B89BCC04E58CA62D <= |I8F57B8D98905C89F4D3B91CA626C25BA ;
I1877CB8174894BB7A9732E91A1794AAA <= 1'b0; I7E04E8229BE60B48AAE3E1EB6511163A <= ID22BB0550BCC1515614C8142FADDA171 ;
I8D181359467F27637239CDAEE8A2F45A <= 1'b0; if (I5FE75BE614D4F52DB327549B36203350 & I0AAD559CF33A5CBA597990658774FEB3
& I923204A95D8CBB206587CF32BEDCF4EF ) begin I7E9516402D6933186513EB5B37336278 <= I3C7A9FA839F554D8898020C4831479E2 ;
IA1EA4D4C05E159614ABC1E6D9CABE3BB <= I74A0936EE8FD1443A2C6745A4F3F6B5E ; end case (I7E04E8229BE60B48AAE3E1EB6511163A )
IAFB2BC0EA796EA2F143B022C32D56FCC : begin casex (I91047088394D6A4116575942899FC337 ) 4'bxxx1 : begin I6B25926923BB34891F18EDE430675796
<= I1A3B3F253A4CAA84340E1092DB0AD78B ; end 4'bxx10 : begin I6B25926923BB34891F18EDE430675796 <= I496D2BA2FDE6A39BB367B7EC043A5D8A ;
end 4'bx100 : begin I6B25926923BB34891F18EDE430675796 <= I0C9CD4F205090AE575352138FEB9E0B5 ; end 4'b1000 : begin
I6B25926923BB34891F18EDE430675796 <= I5898D0798C075683D57F7DA612ED3F03 ; end default : begin I6B25926923BB34891F18EDE430675796
<= I9E0B4C1FB5C57E21C6F98D25B6A3CC40 ; end endcase end IA7E2C061B23F9C2D79751962637FF9F8 : begin ID0A5ECECBEC8CE692F380DDF069E842F
<= {(IBC983AF54FD90EA2AA9E3DD139A3B818 | {5'b0, IE46783A1FBEFC54C8AE5AC3DF183049F }), 24'b0}; I612E93B17FEB6E7AE6FD9448B52CA816
<= 1'b1; end I0FBF38AB1DE3B938794F64EFEB6EEF04 : begin ID0A5ECECBEC8CE692F380DDF069E842F [31:8] <= {I7E9516402D6933186513EB5B37336278 ,
IA1EA4D4C05E159614ABC1E6D9CABE3BB , 3'b0, 8'b0}; case (I6B25926923BB34891F18EDE430675796 ) I1A3B3F253A4CAA84340E1092DB0AD78B
: begin ID0A5ECECBEC8CE692F380DDF069E842F [7:0] <= (ID2E840891AA711130477F703743EDCF7 [0]) ? I476BD51644D400EA02C9B74EB861DDDC
: I961C4AFB4B34DE00139652E84686874B ; ICBC89A2A67F0564ABA5BC46C474021BD [0] <= ID2E840891AA711130477F703743EDCF7 [0];
end I496D2BA2FDE6A39BB367B7EC043A5D8A : begin ID0A5ECECBEC8CE692F380DDF069E842F [7:0] <= (ID2E840891AA711130477F703743EDCF7 [1])
? IDC0F38FB5CB3DE22405E2C1C80579AD8 : I508C4D4DDDB2A017FA853AA88EB418B2 ; ICBC89A2A67F0564ABA5BC46C474021BD [1]
<= ID2E840891AA711130477F703743EDCF7 [1]; end I0C9CD4F205090AE575352138FEB9E0B5 : begin ID0A5ECECBEC8CE692F380DDF069E842F [7:0]
<= (ID2E840891AA711130477F703743EDCF7 [2]) ? I64BD3AC45F8233E09BF36BB23F632819 : I4247280CBF50D75967C778AF3206D432 ;
ICBC89A2A67F0564ABA5BC46C474021BD [2] <= ID2E840891AA711130477F703743EDCF7 [2]; end I5898D0798C075683D57F7DA612ED3F03
: begin ID0A5ECECBEC8CE692F380DDF069E842F [7:0] <= (ID2E840891AA711130477F703743EDCF7 [3]) ? I68321D6CE308BEC2F016764C8A9FCEA8
: I72BD5161F8A297C6D1D0560048EA1612 ; ICBC89A2A67F0564ABA5BC46C474021BD [3] <= ID2E840891AA711130477F703743EDCF7 [3];
end default : begin ID0A5ECECBEC8CE692F380DDF069E842F [7:0] <= (ID2E840891AA711130477F703743EDCF7 [0]) ? I476BD51644D400EA02C9B74EB861DDDC
: I961C4AFB4B34DE00139652E84686874B ; ICBC89A2A67F0564ABA5BC46C474021BD [0] <= ID2E840891AA711130477F703743EDCF7 [0];
end endcase end I2512657214BD8CD9D7C9E46341FB6960 : begin ID0A5ECECBEC8CE692F380DDF069E842F <= 32'b0; end IA4F9276F2E3EF93B14F2B0FF3B2DDE74
: begin I1877CB8174894BB7A9732E91A1794AAA <= 1'b1; end I3AEAA310DC2EB1E6D2E2AB4DD0417BA2 : begin I612E93B17FEB6E7AE6FD9448B52CA816
<= 1'b0; end I9CFCF3FC76F8BCD4AA7E722E67E01A89 : begin ID0A5ECECBEC8CE692F380DDF069E842F <= 32'b0; I8D181359467F27637239CDAEE8A2F45A
<= 1'b1; end IDA65D1282C0B7B2A86436F0450F882A3 : begin I8D181359467F27637239CDAEE8A2F45A <= I8D181359467F27637239CDAEE8A2F45A
& ~I24C403550AE065D7D1B7266142886226 ; end default : begin end endcase end end endmodule 
  module IAC6C4C771C836211892F0FD3F47BC076 #( parameter I857673E5DE2CF777499EE369473CBCCC = "NONE", IA874AED52F9C16F13B580898DA0E85AC
= 0, I45E74A319CD545DA84EE876844F12DF8 = 0, I212658651766EFCF73257AF1E3121AF8 = 1, I2610FF174BEEE098C8D9C9374191F122
= "NONE", IA8729443C3DAFAFDD37A6BED4B24F26C = 0, I08EC85B0527EBF111FDA96E4BD71B6BF = 1, I6C75B7796A1597A63620710B69C04958
= "NONE", I86AD8EB6B8FA8A1AA6EA64DE4357E4EA = 0, I5C0FF6EA47D5544D48B9200C35F2015D = 0, IED6EFA8FE915B71B8E198535343CFBFB
= 1, I98F26EACDFB5625667BCAFBDB2867748 = "NONE", I3CAEAE4A6B7BA30F88F0945373893582 = 0, ICC1064DA289312A92936196EA26F0023
= 1, I78F9B7090517BBEEBC1543199FBA4D34 = "NONE", I731C578B2B8A6173399D3CABA7E98889 = 0, IE18DEDE16538C154B2EFCB2652C25FD5
= 0, IB6EB169241E23C32C11DDDC27322BCE6 = 1, I83476C8D11033DBF952882C55FC0E55B = "NONE", I156838D82D20DC7C269685B24CB4A8B0
= 0, I86134D1B828E3E59B9C4B66EC0920D98 = 1, IC2EB58967FBD1CD5C54491738F4BAD86 = 24'h000000, IBBBF11BAEEC8458B08DFB6E2D9D1C850
= 16'h0000, IA54DA90446D375855AF33292D2570A3C = 0, IAD54DD4DF3ABBB4563A2B75498325CD7 = "INTA", I02756A8C58D5B37B7049B7F6FA2073B7
= 8'h00, I1066D287D755AADD24EE379E400F8DA8 = 16'h0000, IE8C1215A45516D3178A8A93152E05EE2 = "NONE", I6A67F4FE467D33BBE90E5158D72171A4
= 0, I8F998DCDBE9627EA583F7BB408EC780D = 0, I8695C513BA5D9DA307CC481D6AFFB133 = 1, IEE21CD471C5E4E6CE83A164513BC7722
= "NONE", I56DA37D670BDECB81356B81560DC8649 = 0, IB36C0E6BB9CF8D4E4A2F31086369A6EC = 1, I6C4BB963A9FEECAA07E250007DE29E69
= "NONE", I7725F462040C54BFDFC296100F95D5D0 = 0, IC022347DC0BBA44450EA061654CE4130 = 0, I8DFF460C39C720D8E01DF9AD54E62457
= 1, I128970AF889EC52F4195C246A49524BA = "NONE", I61E4D6D4FFCCB1C283902514C76CD3AA = 0, ID0832173F4D69F0B96DB00FA9805F75F
= 1, I171E938E7CDE23987F02EB923184A5C3 = "NONE", I5A509B803B47567D6FA4F4CB4C6AA95D = 0, I2C1FDD71B618A0C398964466A5958BF0
= 0, ICE7C691E1DC04B92371B76DCE234C732 = 1, IA9D9F2D7EEC92A228D6CC71EE9A86E0E = "NONE", I7356A0718B40AEF099CE99273A8CBC19
= 0, I4521B8E3C71C6E5D7639756B81D56C58 = 1, IB52E64F4A5E8239ED2BF949AC0702ACE = 24'h000000, IA5A53C930B674A8F9761966972CFB6F6
= 16'h0000, I97F18A3381F2546EB21E07DF7628912F = 0, I2FCDB5B825200EDE4D7757A0621663E0 = "INTA", IE50492CEE03959C13AD5E521CC7F2FEF
= 0, IC745524098FFC5FBA778DA59D2444D9B = 8'h00, I7507C2B666C444A66EDA2CFDB6DCEEB9 = 16'h0000, I1A39FC80F18CFB225DD25F1158A43FEB
= "NONE", IFA1CC1A50C8D64B9481E806D15AF3CA5 = 0, IF089B8BB6C2663DE1CA53AB4AB67231B = 0, I348F387B0CC3540AF0215535F676D5A2
= 1, I3AB6DCBD252A38D5954C33DB9CFA020B = "NONE", IFE55C92252D5A4FCF3878CC98FCAD612 = 0, IC2181A40E4750EEA118AA81ABB4E415B
= 1, I813CE6D8049DC9123C58691D1DA81B59 = "NONE", I50243AFBCB64F92A3F6EEC157034F4FC = 0, I38E6C6DF2535A2049746702855108B5A
= 0, I0FFEAFBF23F15260885D040F12B66960 = 1, I31E80F0EE05B52A92941F617BDCEF890 = "NONE", I509611AF740C942BA82FB9ECE7BA4E67
= 0, I586C95E6CCC79680B179527AE8977C4E = 1, I39D41D0CFF63339D485BDBCDBC3A8729 = "NONE", IF833CBC3D7A215E6C5635F3F07A09365
= 0, IE106099B16008BAE163236DC5CF4EAFE = 0, IC4C3CD51A29DC2F222334D23407BB4E7 = 1, I7C988FF99F8B28AB1CE2299774306236
= "NONE", I4FF1FE282379DCB83A2AF4F7A12AF6CA = 0, IB5B3486ECA0F911FF5D92A37ECF53B4A = 1, I0B5E80731173820DE30A1D6C548B918B
= 24'h000000, I8A848F283F0A33BC04B5173E5E3FE015 = 16'h0000, I0069A39965C0330678D64B612F60F78D = 0, I30A298A8327798F01C20DDAD6A556FB3
= "INTA", I0B3C14F69FAC563649E26679A3D8B1CD = 0, I4EB1044CFC38A54424DBAA59B9641ED6 = 8'h00, IC920957C9C4BA12361B2EB75CD52EA74
= 16'h0000, IB231E22D146559D11318B25AE0BA8C7A = "NONE", I7377F8B5325C7EE7D12D8B4B6A18183F = 0, I17C1305CE886D24D942A2A62C4DB3617
= 0, ID926607BDA4008824BC8A9A1B67C04B7 = 1, IE4511A2FC6AD3FBAEAADD1EF75F0B773 = "NONE", I0B29563399BE9E04B2FE3DE714C7DCE6
= 0, I698853A251199BE8A5753717E876DA52 = 1, IA3BC4D015F529FD7E88E1370A882D0DF = "NONE", I3463AC2A02018CF2288043A9C3E47A4F
= 0, IFDC235A84B81F7EB6EA5B1ED1F71197F = 0, IF0C0D849F42A4C05A7BF373811D5F5F5 = 1, I59B19D300B55C10DB1B10364E9E59201
= "NONE", IB1CD9FD007D322042A1087AC76B782B4 = 0, I6A959CC2CFE148A0D8579A1CEE0C6699 = 1, I1953E43D30396B1EDBD48DAD13C6A240
= "NONE", IC02B62ACA36F1FEBB031FE435BA48A9A = 0, IAE6C36DBDB6FF8E962D96D8F1FB95CC1 = 0, I82E91D4ACF151209B3234E6F867049F1
= 1, I9806BFEA675277E4572CB4FD0C9C0D8C = "NONE", I802B81175874E1E34C3E4EE6C7F0B969 = 0, I00773A8B25BA28541FF04BC530185E7F
= 1, IB2267C4E34709B9CE9D697340B9DA12F = 24'h000000, I37AC0331E13434E399C90A5408FB09E2 = 16'h0000, IC69BEB80DB094A65F3DFB0265F8616DE
= 0, I6C4A37BD8E4A0A1D9639A3FA64D5F8C3 = "INTA", IFA272F301A5935EE15CB134524665363 = 0, ID969B30E2BD8213873A2D19FFDEF204A
= 8'h00, IC3F1AF003F5E2257563771F88647B5FF = 16'h0000, I21752C34E9BF9458DB0D20BA11A8898B = "NONE", IBFD9199C154D56895B673A496CF82DA3
= 0, I900E9757930519C7865CA2247E6CC23A = 0, IFA7D0D435AE6BBF59445626F82B8B26E = 1, IA794CD2FEB24AB956EC1914852D2E7D5
= "NONE", IAED1399D2D60713A0101069DD427D0A0 = 0, I72E6ED810779933C7E2125FC345DEC0B = 1, I3C7842C10567F9851F14519598E7EE93
= "NONE", I1DE5880AD46DABF7282A3FF245F71602 = 0, I7747208BC7A624CD71D5BB421E9EE4A4 = 0, I4103D81EBFB4946FA8F9593A8B7DE5C8
= 1, I858B464778E6994385995C3205FB37B0 = "NONE", I785E686713BEF380843045D4DB00E51C = 0, IABD30C53E56587015015FE5F556929D7
= 1, IABB4198D13BE4058E856EBC11D8D6565 = "NONE", I0405497FA63FB5AA449F0C813D8E8F89 = 0, I6F86DD61D81AE7AE015C945BA5CF8828
= 0, I69C4352219E15BD98C0B6A7428BAB037 = 1, I68ED8551754B5BAA65EB2F191A697C4B = "NONE", ICE0C22941CF3ECFDB4B47576E4E4A06E
= 0, I262F500CDAF1182E64A895FA5F58D006 = 1, ID88F3DF54AD4CA3D33C94EC1E1B5BB01 = 24'h000000, I8F019158F18BA70FE5953E859D4BA891
= 16'h0000, I4046611EA3EEF60ACE26738C818FDBA2 = 0, I78E815C8C6F11755E08393F339C5E874 = "INTA", IE690B7723F136DA02896C0728DDADB49
= 0, IC377F0EF36016932385B3B0988B91B0F = 8'h00, IBDEA2513680CC11B2E5E42FB17332F70 = 16'h0000, IDC77C35F0E8480627E0F64F68D8A39ED
= "NONE", I110F59F054A1064BFB27909E2370F028 = 0, IED76B05540143124D123636B36A006DA = 0, I96B06C30CEFF410BD39B69C003D2AC2B
= 1, I2050954950618B2F390C43E2A3A4A814 = "NONE", I3F39386711BA6D94D8C7A1C5710875D6 = 0, I3011FF9154FC5D6F394688805C3D9B33
= 1, I08E7BC06415AD0F55BE9EFFEB79B0315 = "NONE", IB069DEA93E56D26CAB0E5B9C9E284CDE = 0, I5F80A9459505144CBBE328F0713782CC
= 0, IC88E0007329C31C00B55FD745AAD6590 = 1, I102247373FC0AC7EA52B3EFB2A5CC280 = "NONE", I750129419895285C7D4ABEB3C2FEEE71
= 0, I2CFDEF4EE4DDBFD88BE646118F3E6FE2 = 1, ID42754EA33A6C985294D5AD602396DA3 = "NONE", I6FBC4AA1ED36E030778F1A24E9C9B2E4
= 0, I15A258E402E001F63FAB5BE8DF569399 = 0, IA2FE22B25B2F0C96B10399B2FB4B7C81 = 1, I36E46FAD7B2BA4DF9270A70F4921CC43
= "NONE", I0500A389ECC6C6D86EA16632126031AD = 0, IFF2CDD869828E984763A775FF1821810 = 1, I4A7FAB30233B5A9954B6B6AD08DCADAA
= 24'h000000, IC7B583F6D8F8A6C3C62D45FA87D50A19 = 16'h0000, IAE03DAE231BA40E8DD1C02D38068EF8A = 0, IB842E33563B3EE1795267FE015C7B1A0
= "INTA", I55BE27080C370AF723A4FE096014E875 = 0, I229F764F8E53B82969E0B6B9234098CF = 8'h00, IA9807BAB69B1AFAF9739BF86D99A92C3
= 16'h0000, IF02D8DF664D45B9699745A4C477F4220 = "NONE", I553DE26948BD8999C232161660D3E8AF = 0, IB99020DD53AEEF55E5DA5BF15890E9A5
= 0, I0108C021E74AB8DE1357A170111B08CF = 1, IDED06CF1ED1692C601F91B904599696F = "NONE", I7926E122D54A321BCD3309E19D9A0183
= 0, I48C74401BD4D3F04619117E263213AFA = 1, I40F4EF6A18605258D6F6893B593AA318 = "NONE", IAB56F2CB5ED41158B5A0ABE2FD915084
= 0, I11F59D9A3377C9C28FB84219B4A4E4DC = 0, I3BE4D977225B6255BC284FA193DD9241 = 1, I6A49481E89496C888774F840785C0BA4
= "NONE", IE19B87A06C26E07981B4C116F5E878F7 = 0, IF587F6E4A635FC1DA01C698D24B80510 = 1, IBF68DF087726DF134221B625725579B8
= "NONE", I9F10A6A60E1AEDF0BC22B2ED2686E4C2 = 0, I10394C1F82392903C22C104CEC600C4E = 0, IE4A74A61CDC56044C199B3C3D606B08E
= 1, ICE73FC6522779AED50B02BB41E81D717 = "NONE", I25D595F391F999FD69AB7E7B5B1FA99C = 0, IAE37CBAA4815C82EA96E8FA0802F7443
= 1, I50BD52F5094656ECEC3714E0BAE6B0DA = 24'h000000, IC781EE34DC62D08174F1793A9E3131B5 = 16'h0000, I7568F6D9A53738CCE095CE231BAB3F85
= 0, ID23C9147B8CA6684051791F38B473984 = "INTA", IB2560D175E4507798B84D6E659FD6373 = 0, ID873CC05798FE57AF43DD3C4E138769B
= 8'h00, I70E83CF258ED794C3E9EDE1260BF5578 = 16'h0000, IFB72ECF29D30B02049C030502F330CE7 = "NONE", I7E6B00724A48BA5DD1C5E397542EDDC2
= 0, I5C146FC803FDD1163A6BAEA53E6C5468 = 0, IE3404D24C7B1FA263F2EACB5CC85BFF6 = 1, IB23260A86DA99A28163B5E233CA42605
= "NONE", IEF68A43ED89112E53191106DBA0EF113 = 0, I95CE19A3BB94C8A24A8E3F3482EF6425 = 1, I7A84A5F1499409083F731D2A584D2D42
= "NONE", I76069160333C4C8E92944FC3A3827ED6 = 0, I8EF5BB87B22B910665D13A80C6724D14 = 0, IFA5339CE0FEDFF3B45CF3C0167564EA1
= 1, ID3A400426A266A6F4E75F7686B9028CD = "NONE", I071A2CF414FF8A814D779E1F54247BF1 = 0, I3F7B58F167F56FB985F8908CA1B7E3AE
= 1, I62A26688D23065F69E9B9D6339AA01A5 = "NONE", IE4774E19FB83A84DBF540368C45EA3A3 = 0, I5ACFA0E62CCC520EE4DA1BA399F1B7E6
= 0, IF1CB2B99D8669C68B68BC468C83323DF = 1, I245B45EC852C565EDD1AAC06E80DABD2 = "NONE", I59DF7AA363A19A361E3A844AD6039C40
= 0, IAF2433492FE33171692143422229D319 = 1, I721D73CBB11DB0EC9DF361993F6A92EA = 24'h000000, IE0DA0C810288CC00DF1F3AE622FFB08F
= 16'h0000, IEB4CAA0AE4F26FAC1DAA6B9884179DEA = 0, I070D33CDFCF15FB7B4DD88019C0E39E2 = "INTA", I25B649490B20A1FEC9A1AA60AB0C6D5E
= 0, I8302D4B9F46621BBB824B1CC96E2E724 = 8'h00, I26BFDE09E6F548FBAC63338567411C7E = 16'h0000, I46C5269B9FB24EF04CE2CC341C288EC7
= 16'h0000, I3C9AD458B89B2FAABD743BF4E13BF421 = 16'h0000, IAB32DAC10CBDBE04FD5EDBF7A576CAF9 = 512, I394B9366718FFFBF01944193881668C1
= 0, I66C185998F46A7148163982E39BCD296 = "ECP3" ) ( input wire ICCFB0F435B37370076102F325BC08D20 , input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 ,
input wire [63:0] I8B1798242C3B0E655181D0D365813614 , input wire IE145222FDBDC80109E12FA72D3D3C655 , input wire
ID43AC1009727D128F1C5DFE4640CA5AB , input wire IB610431939CB8180EAC2403672BAF58D , input wire [31:0] IEE7B9D1B054F5CACBC10351FC32D7BFA ,
input wire [31:0] IFE8155182FD754C22D6F7FDA1F1C1174 , input wire [31:0] ICFA3AEC9D2E8697060447D8D8EB18A80 , input
wire [31:0] I81D61D198832883CFD88EB5DEB88A32B , input wire [31:0] I1F5A786F105B576AC15A6F25EBFB89B8 , input wire
[31:0] IB9B532CA44CE4054811AB748EDD0922D , input wire [31:0] I7FE73B332A2A7E273F8EC82CC2A0A9D1 , input wire [31:0]
I8C784B1A25E6B5F5402709647F921D20 , input wire [31:0] IAFB7D4809B407BA0A70ABF120DF37844 , input wire [31:0] IA69AD6BF563BE83DB737C644B2992470 ,
input wire [31:0] IBBC01C0CF0EE486327FBEB391C90772B , input wire [31:0] I147607D1A744B7E8E0F3050C499F3A23 , input
wire [31:0] IAA6C398FE19CA194DA9436764C94079A , input wire [31:0] I6375C05D4E0F58631C8731FD2B26A7F6 , input wire
[31:0] ID25293C6DC5461B1A3E61F7A7614A6D8 , input wire [31:0] I7E0B227F296E6A7FA770C68AB70324DD , input wire [31:0]
I1187CE134A1A3347BF94366BE4D44B3F , input wire [31:0] I0C7C3FDEC159F63C155144A19841E5BC , input wire [31:0] IF0C365E1D4BC8B2941DE257EF66C8FE4 ,
input wire [31:0] I1646E818A90159BC4FF7AA119272C460 , input wire [31:0] I05AD49E3884F0E62FA36DCFB88E5C22E , input
wire [31:0] I348CE8EA5A014339F820FDCAFC214867 , input wire [31:0] ICF2AC2986B60A3FD41ECFB74C4756D10 , input wire
[31:0] I13B899B342E8552CACED9E20E0F5FD83 , input wire [31:0] I068B3206EC02BBE1225E3FD649DCAC3E , input wire [31:0]
I15D8A1D8934ABE732F753BC8A130129E , input wire [31:0] IFE8F569C18FBA7444D4832F2CB5D2D69 , input wire [31:0] I51FF9F99E3F92A151FD3D6BBAAC89FB6 ,
input wire [31:0] IA4118298EF0A9C92D5D3ECB07C8AE533 , input wire [31:0] I7D032A1E448C6F22898894E594BF2DD3 , input
wire [31:0] I67444F97CA6B95448FAFAE30BC1EA4A3 , input wire [31:0] ID449FF330193AAA4C7942F23F18CEF54 , input wire
[31:0] I3CABF30E4ECE3E02DF7BB2FAE8895026 , input wire [31:0] I46EAD98AAF05965858087C6CCDFEAFFD , input wire [31:0]
I1967BD95F38270D97B0A4B182C5D8F0E , input wire [31:0] ICDB8224D569BB5A5B320A26E2B451BAC , input wire [31:0] I8220BA29B6C07A3A107C2B3234F5FB06 ,
input wire [31:0] I7DA2457F5006629E45D78C4FC855DCF8 , input wire [31:0] IBB764C0D62FD349F6FB3F52A8C78424E , input
wire [31:0] IE074E5B8DF895724AB3B5023BAC298BC , input wire [31:0] IDA2FA24095F53E4EBBAC1E30772082B4 , input wire
[31:0] I27FBA72EC841BBBDD25E028A08A3F06C , input wire [31:0] I4FB68E387DB515A46DAA2DABF6E0D1D8 , input wire [31:0]
IBA4DC2E68E546946B55995DB900F74F7 , input wire [31:0] I28A9F4DDE0D0FFADF8668EFA99C6DA03 , input wire [31:0] IE02A2D602D1C83798270DD49EF6A4D23 ,
input wire [31:0] I4DBB86A2215D89E37CDE4EC7DC8435C5 , input wire [31:0] I8DCB72E575B62CC266039827C0238E34 , input
wire [7:0] I3C7A9FA839F554D8898020C4831479E2 , input wire [4:0] I74A0936EE8FD1443A2C6745A4F3F6B5E , input wire [2:0]
I369BA2FFB5D41DF25F9BC3AB126D6607 , input wire [IEB4CAA0AE4F26FAC1DAA6B9884179DEA + I7568F6D9A53738CCE095CE231BAB3F85
+ IAE03DAE231BA40E8DD1C02D38068EF8A + I4046611EA3EEF60ACE26738C818FDBA2 + IC69BEB80DB094A65F3DFB0265F8616DE + I0069A39965C0330678D64B612F60F78D
+ I97F18A3381F2546EB21E07DF7628912F + IA54DA90446D375855AF33292D2570A3C - 1:0] I1C0271AD5E8E9E9164909E468AD0B212 ,
input wire [7:0] I6EC1BE4B18EC6AA3D88A5D45B614565E , input wire [8:0] IB907C2624CE144BCE5A772623C46F678 , input
wire [$clog2(IAB32DAC10CBDBE04FD5EDBF7A576CAF9 + 1) - 1:0] I3FF97406B3ED373B267711109A980AF9 , input wire I24C403550AE065D7D1B7266142886226 ,
input wire [14:0] I438B8BD876741F9B46EB770E92F808B7 , input wire I5FE75BE614D4F52DB327549B36203350 , input wire
[31:0] I3D6C771D05CA1A769E61302C086494B8 , input wire [3:0] I357B3043EDACE3EBECE8F54D79B9F90A , input wire I0AAD559CF33A5CBA597990658774FEB3 ,
input wire I923204A95D8CBB206587CF32BEDCF4EF , output wire [7:0] ICF9D8FD31DFC7D20DAF939C6D75F1518 , output wire
I20CD33DEFBDF51E2A5352736B083738D , output wire [7:0] IDF550B17734BF16B7E410B19BB31E276 , output wire I8ED9B9C1D9F58C5D06A9443AD901E8C6 ,
output wire IA976D63BEECA80DCE31365CF56EC0248 , output wire I5E3CE5AF5C34D232BFB139B63D9912B4 , output wire IBEF3E5F9395E2C7822AE03D6461DEBBB ,
output wire I7E6CFD6A7DCAB9CD2188D044C7D716A6 , output wire I3A34691662384260F0524DD7F650E75A , output wire [7:0]
IC2F58AB5028C1D2C53C6EF47A4975D0A , output wire [2:0] I112E0A79129A8BC6DD4C13647C31F8A0 , output wire [7:0] ID3E7F4B58943229FEE6313A36B3F8693 ,
output wire [4:0] I1FDEC1735547330C00A0B8DFE1FB10C3 , output wire [2:0] IBD6A65D48B4A68CA0D2A82F79053757B , output
wire [2:0] I42A419EB6EB8D11234AC3B2BCA0AE593 , output wire [2:0] IA41AC3CC6BC050DDC172724AB311315B , output wire
[7:0] I31CF69FF368B36B4D6612DF16B3ABC6B , output wire I439AF6D496491F5F7C23217209B43C31 , output wire [31:0] IFE4A8CBA73734C6F0F0A078027E053D4 ,
output wire ID7A2A8B1E9D92B60194D5FAFAAB15208 , output wire IF274FAF97F5BACD693913BB418717A9D , output wire I270ED686C2EF2C1C8B5B55EC4A5AAE84 ,
output wire ID5CCD4858CB5CC1B2EDEC682C7DE5AAD , output wire [31:0] I7D901091F9E0741061C75B54467D48A0 );  localparam
IB26EBF559CA483EACBAD1BCA4C580AF2 = IE50492CEE03959C13AD5E521CC7F2FEF || I0B3C14F69FAC563649E26679A3D8B1CD || IFA272F301A5935EE15CB134524665363
|| IE690B7723F136DA02896C0728DDADB49 || I55BE27080C370AF723A4FE096014E875 || IB2560D175E4507798B84D6E659FD6373 ||
I25B649490B20A1FEC9A1AA60AB0C6D5E ; localparam IE3D0FF95EEFE7CF51F7D6968D26EAB4A = 9;  wire [7:0] I74CF4D6FE5B30BB30E40AFCA2A08A220 ;
wire I60003168A46706B958CCEC72E50AC23E ; wire I111827C337F00C09A8C61C3DCE514338 ; wire ICF847A44ADAE70C9998962202A23AB4E ;
wire IC4C35B8C650EEF422BEF8C68B5A9359D ; wire IB624795CEFFC2094E111CAD5578DAE1C ; wire IB56580C539321C40E6B44EB394A9EECF ;
wire [7:0] I400149787F2546E3D0331041FB8123FC ; wire [2:0] I97E631353C4C7709CF07D5FC5800DDBC ; wire [31:0] I97B15B5DA5A0868F11CDF3929B25044E ;
wire [31:0] I16A1A5B65742A57E7143E981BF286F99 ; wire [31:0] IB4CA57E47B085EE5925036D5223A4598 ; wire [31:0] I2F92739468FA7128C93936C8511AA228 ;
wire [31:0] I25DCCEF37BE2FCC042C00B81ABCA449F ; wire [31:0] I19381BD04F07A020B45A7EFE952EBD90 ; wire [31:0] ID54A2FD9EE0AEAC4E7AC2A4D30D28B9B ;
wire [31:0] IA5469486BB0530B9AA1B819A3C7A9583 ; wire [7:0] IACF97B89AE62537A26788BDFCE846ED1 ; wire [7:0] I01D4C6B20466D26621C6DA5816817455 ;
wire [7:0] I46A701488EBE724B47736C3C7A47A876 ; wire [7:0] IFE63F76C2A46B87271596BE8D0FFD21A ; wire [7:0] I21EE6CA5EBC86B66AC5EE8AF763FB838 ;
wire [IE3D0FF95EEFE7CF51F7D6968D26EAB4A - 1:0] I56519DD369C66F1A0EA1EE3D2398E0EF ; wire [IE3D0FF95EEFE7CF51F7D6968D26EAB4A
- 1:0] IC0667A37FE3E5F8D3579C6AEF86F5C24 ; wire [31:0] IED75BA58ED5F09B80AEBB5C4531DD96E ; wire I86E103F0E5684240BF4D6AD4E9635C7A ;
wire I6618736D0C53F4C6D20F8C252BF264AD ; wire I5917F25EB5F020E0FEEB03EB956B3110 ; wire I9818F0A46507B01B5AAD29ECB3D36F81 ;
wire I0EB153824311AB3255F80A6B20F59828 ; wire I6A77961ADE4327F78C7D008C5DA7D184 ; wire I8C1666B519246534E1C4722652FD1823 ;
wire I95628D4658FCAB1EADD1EBA1F6294ED6 ; wire I841AB9A2043753D035FC3A85DEFAF1D2 ; wire I711EA37894AB982C997C1497E71677B4 ;
wire [2:0] I42DFCF8044FC66463EFBDCD6F2C69AEE ; wire [2:0] I999118EB4E0839ECF8CF049C93027B49 ; wire [2:0] I6080D873E932E26F13608A1D73FAE7C0 ;
wire [31:0] I1179A173C6F4C43BA9C3B71086E48486 ; wire IC99E8E0D5BAC180B4FAC3C67D1618142 ; wire I1C08DD68F49BF5FFE04D852950D9A932 ;
wire I6AF9911F8AAC2F653011D5D8ACE5F433 ; wire [10:0] I7D2B5C97BC25D475F870C1BE7E21B697 ; wire IF082298B35C4A83318C3597AC50DA20E ;
wire I762EB11F447E9FE5C306D10B1D44F3D1 ; wire I7ED71D3164ABC636AC5046B7E263FD03 ; wire [31:0] I6795B29551221467FFA6B7172DDA857D ;
wire I25D510B1A7EEBD7D688C48A4050B0A28 ; wire I85BF4AD7C60BEA5045D19571D851C992 ; wire IBF1BA20BCDFE79989AD3C8104A1024A4 ;
wire I4B2CDC61C9F80778CDBA134570DB93A1 ; wire IB3122CB8FBD2C123E9D9BD0599AE41D0 ; wire I2A46DB8D4D31FAC435A47D582BA0E704 ;
wire IF6683BD4A4C0331D12A89BC5CD3FDAA2 ; wire I40DCE993F9A1E526661825B1281A7DCB ; wire [2:0] I9A3A1B70A9C668CF11493348B519FF4B ;
wire [2:0] I09A93891DA1B4315581C9B6775306EC6 ; wire [2:0] IA60C7697AAB3A707DC265C02AA59526E ; wire [31:0] I3E4C4B769B824746306BEC19D75E1A23 ;
wire IA2B524351B6A8AB3A2FA7E1B456ABE67 ; wire I037B294714AE918C1D513F83470C0190 ; wire I6FE2694F3F3B5838177CEF5992A016F2 ;
wire [10:0] I976ABC47C39290CF3E29B8773D338ECE ; wire I42864A73C6A7A061BF0E25880AF8AE9C ; wire I24FB1AC5C4A1C96F7DF559EABAD558C5 ;
wire ICA544D75FD0BAE421ECEFDBC4207F6C1 ; wire [31:0] IEC017B3AB9F16AE871D5253A5257D941 ; wire IB1AAAED8469CADFA3AB4BF806A8466B6 ;
wire IA6774F4F4F3AF83C6A9E233DB00F89A0 ; wire IFFF50035216FD68A74F8164F0EE74689 ; wire IF9A16909C25386742335A246DEDE12E8 ;
wire I5078F81AE0F5DCD4CC2ABEE2CEF9C827 ; wire IB55475954FE95F83F22B1C2FB76FAEC7 ; wire I31980ABC07D19BA89784085C7754DE42 ;
wire IE1F9397E899B4E938A0D54FC51445C13 ; wire [2:0] IDE0F2D42601304C0E0CCD60778B3938F ; wire [2:0] IAF2A92B584FD036A9F751EB8F3FA7ACD ;
wire [2:0] I5CF35907FA895D81AAC1AAFED86DBE1F ; wire [31:0] IFFB9EED620356BDFB94697DB3606174F ; wire I2C072E656BFCADF4877B42244D6D2307 ;
wire IB96A9322FAF5941DF70737CA69F152A3 ; wire I5B92AFCE2F6F881BA10FA726B18BB692 ; wire [10:0] I60F6B756CD1062B40CC02E1438F28711 ;
wire I746F8C8440813F740701D80A6F08674F ; wire I9625E96E33563830A2A0ED7263124B10 ; wire I1B43D1CE930FCA067FA31726F2C15FEE ;
wire [31:0] I697639B04C0F4B6F9764F8122329FB7C ; wire I1E1A1AD224EE52C02213B0661856A826 ; wire IDBF2DE7607B69A821EF14BD65A75A2DC ;
wire IB35E0CDEF8AAA93EF9B0047DE75BCDB1 ; wire IC5663A92559813188629C72D2AF75E2B ; wire IB7ADE2C78FA2211545637C290CFB45CB ;
wire I38BDB4EBCC779338E7AF863601C4853E ; wire ICD34F2C7357A369358E7CFBC3D425106 ; wire I081CFEF0428EFE96BD06A8F2EE9DC2CD ;
wire [2:0] ID34187ADCB71E296DE727A7573E76A15 ; wire [2:0] I5B6B84BEB62496031A951D18F8043152 ; wire [2:0] IC21D6CA5169E489082288A960FB9DDFE ;
wire [31:0] I0D8A716B0016AFE64E7F7977A80A253A ; wire IAEFBAA4728FB6854C056C8E4C0691B3D ; wire I1DC328E1B03775141AFCFBB60C78CDC0 ;
wire I3ABE7E8A0A3ADCF18D9C06A84D938210 ; wire [10:0] I6DA6F40C5003D56BA074AD254DFE4B48 ; wire I55D773F0648256E2B67F14A58A7AE480 ;
wire I0F56078C1F80B8234A46BCE05F251A14 ; wire IA37321C9DB7C6279A1BBB82432DD22B2 ; wire [31:0] I3C0E217327A8665923FDC969639C89C7 ;
wire I22F7EBEFD72C22C64DB546CE211C3C33 ; wire I7DA4C0DA5661A2191D932C4F426DE5F4 ; wire I17B065631E7403BD94AABA998687E920 ;
wire I2D58D8090233025B63B11977CCF7A6FB ; wire I79527CA6375BFC9B46B48DEFE32DEEAA ; wire I270710745C28824E285C2E05FB618D27 ;
wire I765A5C6CB6D2AE7496EF2BE962529E09 ; wire I9C559D18449178998B7475813A7D0CBB ; wire [2:0] I7B62DE436B5B4C0A20CC4FE1E5D6F91D ;
wire [2:0] I56408FACA355983EAB06294FBFDA5C73 ; wire [2:0] IDAF814B27DE872458FE905492366EC1F ; wire [31:0] I88DEF602C28E2AE7FCFC75761E9DF8F6 ;
wire I6434FE6B1DB9B4DCDB82F1E568D8A5AD ; wire IF76FEAB2FA7E91BC33928D6B232B6040 ; wire IA3A543EBA3F35D293D9F9A372241FFB7 ;
wire [10:0] I6913053E317EA8A5066057EFF8119A7D ; wire I96F424D83A110B76A1E3957956BB0EEA ; wire ID24D46A573CB38B617C5B4569142A8C0 ;
wire I097D8CB350937ECACE8C02CAB12CF7F5 ; wire [31:0] ID04E1BCD61D6D921C4E551FD2CE92041 ; wire I0ED491A5B7F42029CCB818A7A566A126 ;
wire I64422991E0FA499CEA26156FB729091E ; wire I1C44B39C210FB0191DFBF4FF9B4EB5AC ; wire IC3DC126AC872E9080FFE257241E00572 ;
wire IBCCBF2F5A49A76D461A7479DA2813EA7 ; wire IFFE90484B4E519D0DD55AFC0D9379B2A ; wire I6FDDB4608592CC601F82E29CF03F58E2 ;
wire IE6E0B2D716FF39D4E07D15E9EAAB04FC ; wire [2:0] IA2F68AF483F09457F392B22939441F47 ; wire [2:0] I8238B208D31228316827652162FA0720 ;
wire [2:0] I28192CB07D936DD6F915E872C9D77566 ; wire [31:0] I98308209671212A3C88A9644B503FA02 ; wire IB4C822D6BFAE40F12254437B18142B8A ;
wire I30157CAB406F288B630EF42C05ACC134 ; wire I82635882370B55739EA7454635CE3A41 ; wire [10:0] IE38989B54E8F0643FD2DC5F4F7B5BCC6 ;
wire I42E863B8B97EAE3620723BFD560E96F6 ; wire I5ADEE764CD8A8EACE17ED8F55EC633AC ; wire I977D818DD621CC225F1001F838F63684 ;
wire [31:0] I56C985EEB74E064645781DE4618A62B0 ; wire IB9FE9C794CFE66C9E361CA5E0C2E0ED0 ; wire I200264A7B4F7EBBCB0636F8B0C705433 ;
wire I5FCD09AF69B4D4969F86A3686036D558 ; wire IECF63199E2CFF774FC2362604C428EEF ; wire IABDBB85ACD3277D447B4FD8665EA150B ;
wire IB77F87CED77CEC2F6256375F35443CD0 ; wire IAF3303768435E5C76A60A5987AF1CD0A ; wire I2130A737A8CF0DAA0688CD61C692C53A ;
wire [2:0] I009BA1F74DBCC8E4177F1254D60DCAE9 ; wire [2:0] I3710541DAEAC21250982ECECA6E16679 ; wire [2:0] IEF2F499EA80B8075F4C485F59E3AA64D ;
wire [31:0] I386D96EE2FCEC8374B24F3017B94BD4D ; wire I11E1C086CA3C13B481A5977B8AD8694F ; wire I5C58E3085FDB240D9A5DD64A9CD3A30B ;
wire IE0683883BF201CF74ADDEE61816AAD96 ; wire [10:0] IF4776D1E9086F7D152D43C91A22BC985 ; wire I176659D1476D3660538A1C22EFD75A83 ;
wire ID0B88392A9310E618D259D3AE74555DF ; wire I2467937CC723EBC133B60C885A06C7A8 ; wire [31:0] I3FC95340E6F01F64D548828DC3B2A0FE ;
wire IDEEB7827D919A8134F28A8BCC126AD5D ; wire IA7846F08DDB80EC63AA4A9EC1770A3F0 ; wire I93A8E9B4C6DB1D603A05A9591C4339C9 ;
wire I17CB952AA0F6F5C6792E1381BEB60CA3 ; wire IEB1DC53BA14A2028F346A4C10651DA08 ; wire I7616B3B0828958A3CA36203B840CF4D6 ;
wire I246B1D75EEA1239D65C20304AF791CB4 ; wire IBCEA86C0BDF1E124E6697E40D620DD0A ; wire [2:0] I11D20DB2F186022215040429BE705A72 ;
wire [2:0] I73B39CB9A73EAB03AD04B21F62F95224 ; wire [2:0] I700C2FF696E95E1F0C6E6B8EB54971BC ; wire [31:0] I49850943EA73C8BE46401A2FC9B67D74 ;
wire I14F6DF0BCAC12F6EBAD7145BDD4B2D26 ; wire IB85FB30E34AF0B105FD21BBBB73605EA ; wire IE67F175E6F2CC66DDCAD62CCD21F3551 ;
wire [10:0] I58A4869C5AA5FC57B207E7883C179856 ; wire I9DD533FE3D53A79078BF27CC1058785B ; wire I4D0BD33FE293DDEE3A568B64EE8F63F1 ;
wire I42FFAA9F6065323EF66FBE15FAE57258 ; wire [31:0] IE8EF8CF3D14B7C15DC96E6E2DC4BA14A ; wire I18AB4B503F92B00D610DFDE3078A4B8F ;
wire IAF7DC8691D3941B7E52C532F1E8C7FE1 ; wire IBFA78112A3EFE7AB665D3E3A9A588B1D ; wire I94288AE7E6EFEA1989E284E9B2867097 ;
wire IDEB44FD98C3E74E285A47A4BD69A7619 ; wire I3A3A0FDF754EB1C6D50FABC25DBFC696 ; wire [7:0] ICCD7B28178C3803739C5C1C758B836E2 ;
wire [7:0] IC7DB18773990D347CEF55E672D6B2C05 ; wire [4:0] I39A06B46F4E1C11EE4BFB781E3B4F32A ; wire IA513FFA7CDD6BF8E65B629CB494239A4 ;
wire [31:0] I6DFBACFF2E5A466B93A00001848429F7 ; wire I7CA41EFBA3D0548B989711570EA40B95 ; wire IC30C68A9857DD63CE5A51E5943CEB3AF ;
wire I8824AFA21C1B61513D8DE94591B948FB ; wire IB5292E1DAB3B0E7E62E43F792E80D8F1 ; wire ID4282AD4BEFA96986B17E55149DF417C ;
wire [IE3D0FF95EEFE7CF51F7D6968D26EAB4A - 1:0] I81BF37FCB51B492DCA857F28ABD8D76E ; genvar I24501E622BFA6932719D2F78F75F6270 ;
 assign IDF550B17734BF16B7E410B19BB31E276 = {IDEEB7827D919A8134F28A8BCC126AD5D , IB9FE9C794CFE66C9E361CA5E0C2E0ED0 ,
I0ED491A5B7F42029CCB818A7A566A126 , I22F7EBEFD72C22C64DB546CE211C3C33 , I1E1A1AD224EE52C02213B0661856A826 , IB1AAAED8469CADFA3AB4BF806A8466B6 ,
I25D510B1A7EEBD7D688C48A4050B0A28 , I5917F25EB5F020E0FEEB03EB956B3110 , I5917F25EB5F020E0FEEB03EB956B3110 }; assign
I8ED9B9C1D9F58C5D06A9443AD901E8C6 = I18AB4B503F92B00D610DFDE3078A4B8F ; assign IA976D63BEECA80DCE31365CF56EC0248
= IAF7DC8691D3941B7E52C532F1E8C7FE1 ; assign I5E3CE5AF5C34D232BFB139B63D9912B4 = IBFA78112A3EFE7AB665D3E3A9A588B1D ;
assign IBEF3E5F9395E2C7822AE03D6461DEBBB = I94288AE7E6EFEA1989E284E9B2867097 ; assign I7E6CFD6A7DCAB9CD2188D044C7D716A6
= IDEB44FD98C3E74E285A47A4BD69A7619 ; assign I3A34691662384260F0524DD7F650E75A = I3A3A0FDF754EB1C6D50FABC25DBFC696 ;
assign IC2F58AB5028C1D2C53C6EF47A4975D0A = ICCD7B28178C3803739C5C1C758B836E2 ; assign I112E0A79129A8BC6DD4C13647C31F8A0
= I97E631353C4C7709CF07D5FC5800DDBC ; assign ID3E7F4B58943229FEE6313A36B3F8693 = IC7DB18773990D347CEF55E672D6B2C05 ;
assign I1FDEC1735547330C00A0B8DFE1FB10C3 = I39A06B46F4E1C11EE4BFB781E3B4F32A ; assign IBD6A65D48B4A68CA0D2A82F79053757B
= I97E631353C4C7709CF07D5FC5800DDBC ; assign I42A419EB6EB8D11234AC3B2BCA0AE593 = I999118EB4E0839ECF8CF049C93027B49
| I09A93891DA1B4315581C9B6775306EC6 | IAF2A92B584FD036A9F751EB8F3FA7ACD | I5B6B84BEB62496031A951D18F8043152 | I56408FACA355983EAB06294FBFDA5C73
| I8238B208D31228316827652162FA0720 | I3710541DAEAC21250982ECECA6E16679 | I73B39CB9A73EAB03AD04B21F62F95224 ; assign
IA41AC3CC6BC050DDC172724AB311315B = I6080D873E932E26F13608A1D73FAE7C0 | IA60C7697AAB3A707DC265C02AA59526E | I5CF35907FA895D81AAC1AAFED86DBE1F
| IC21D6CA5169E489082288A960FB9DDFE | IDAF814B27DE872458FE905492366EC1F | I28192CB07D936DD6F915E872C9D77566 | IEF2F499EA80B8075F4C485F59E3AA64D
| I700C2FF696E95E1F0C6E6B8EB54971BC ; assign I31CF69FF368B36B4D6612DF16B3ABC6B = I21EE6CA5EBC86B66AC5EE8AF763FB838 ;
assign I439AF6D496491F5F7C23217209B43C31 = IA513FFA7CDD6BF8E65B629CB494239A4 ; assign IFE4A8CBA73734C6F0F0A078027E053D4
= IED75BA58ED5F09B80AEBB5C4531DD96E ; assign ID7A2A8B1E9D92B60194D5FAFAAB15208 = I86E103F0E5684240BF4D6AD4E9635C7A ;
assign IF274FAF97F5BACD693913BB418717A9D = I6618736D0C53F4C6D20F8C252BF264AD ; assign I270ED686C2EF2C1C8B5B55EC4A5AAE84
= I762EB11F447E9FE5C306D10B1D44F3D1 | I24FB1AC5C4A1C96F7DF559EABAD558C5 | I9625E96E33563830A2A0ED7263124B10 | I0F56078C1F80B8234A46BCE05F251A14
| ID24D46A573CB38B617C5B4569142A8C0 | I5ADEE764CD8A8EACE17ED8F55EC633AC | ID0B88392A9310E618D259D3AE74555DF | I4D0BD33FE293DDEE3A568B64EE8F63F1
| ID4282AD4BEFA96986B17E55149DF417C ; assign ID5CCD4858CB5CC1B2EDEC682C7DE5AAD = I7ED71D3164ABC636AC5046B7E263FD03
| ICA544D75FD0BAE421ECEFDBC4207F6C1 | I1B43D1CE930FCA067FA31726F2C15FEE | IA37321C9DB7C6279A1BBB82432DD22B2 | I097D8CB350937ECACE8C02CAB12CF7F5
| I977D818DD621CC225F1001F838F63684 | I2467937CC723EBC133B60C885A06C7A8 | I42FFAA9F6065323EF66FBE15FAE57258 ; assign
I7D901091F9E0741061C75B54467D48A0 = I6795B29551221467FFA6B7172DDA857D | IEC017B3AB9F16AE871D5253A5257D941 | I697639B04C0F4B6F9764F8122329FB7C
| I3C0E217327A8665923FDC969639C89C7 | ID04E1BCD61D6D921C4E551FD2CE92041 | I56C985EEB74E064645781DE4618A62B0 | I3FC95340E6F01F64D548828DC3B2A0FE
| IE8EF8CF3D14B7C15DC96E6E2DC4BA14A ;  assign I74CF4D6FE5B30BB30E40AFCA2A08A220 = {((I438B8BD876741F9B46EB770E92F808B7 [14:12]
== 3'b111) ? I5FE75BE614D4F52DB327549B36203350 : 1'b0), ((I438B8BD876741F9B46EB770E92F808B7 [14:12] == 3'b110) ?
I5FE75BE614D4F52DB327549B36203350 : 1'b0), ((I438B8BD876741F9B46EB770E92F808B7 [14:12] == 3'b101) ? I5FE75BE614D4F52DB327549B36203350
: 1'b0), ((I438B8BD876741F9B46EB770E92F808B7 [14:12] == 3'b100) ? I5FE75BE614D4F52DB327549B36203350 : 1'b0), ((I438B8BD876741F9B46EB770E92F808B7 [14:12]
== 3'b011) ? I5FE75BE614D4F52DB327549B36203350 : 1'b0), ((I438B8BD876741F9B46EB770E92F808B7 [14:12] == 3'b010) ?
I5FE75BE614D4F52DB327549B36203350 : 1'b0), ((I438B8BD876741F9B46EB770E92F808B7 [14:12] == 3'b001) ? I5FE75BE614D4F52DB327549B36203350
: 1'b0), ((I438B8BD876741F9B46EB770E92F808B7 [14:12] == 3'b000) ? I5FE75BE614D4F52DB327549B36203350 : 1'b0)}; assign
I60003168A46706B958CCEC72E50AC23E = I9818F0A46507B01B5AAD29ECB3D36F81 | I85BF4AD7C60BEA5045D19571D851C992 | IA6774F4F4F3AF83C6A9E233DB00F89A0
| IDBF2DE7607B69A821EF14BD65A75A2DC | I7DA4C0DA5661A2191D932C4F426DE5F4 | I64422991E0FA499CEA26156FB729091E | I200264A7B4F7EBBCB0636F8B0C705433
| IA7846F08DDB80EC63AA4A9EC1770A3F0 ; assign I111827C337F00C09A8C61C3DCE514338 = I0EB153824311AB3255F80A6B20F59828
| IBF1BA20BCDFE79989AD3C8104A1024A4 | IFFF50035216FD68A74F8164F0EE74689 | IB35E0CDEF8AAA93EF9B0047DE75BCDB1 | I17B065631E7403BD94AABA998687E920
| I1C44B39C210FB0191DFBF4FF9B4EB5AC | I5FCD09AF69B4D4969F86A3686036D558 | I93A8E9B4C6DB1D603A05A9591C4339C9 ; assign
ICF847A44ADAE70C9998962202A23AB4E = I6A77961ADE4327F78C7D008C5DA7D184 | I4B2CDC61C9F80778CDBA134570DB93A1 | IF9A16909C25386742335A246DEDE12E8
| IC5663A92559813188629C72D2AF75E2B | I2D58D8090233025B63B11977CCF7A6FB | IC3DC126AC872E9080FFE257241E00572 | IECF63199E2CFF774FC2362604C428EEF
| I17CB952AA0F6F5C6792E1381BEB60CA3 ; assign IC4C35B8C650EEF422BEF8C68B5A9359D = I8C1666B519246534E1C4722652FD1823
| IB3122CB8FBD2C123E9D9BD0599AE41D0 | I5078F81AE0F5DCD4CC2ABEE2CEF9C827 | IB7ADE2C78FA2211545637C290CFB45CB | I79527CA6375BFC9B46B48DEFE32DEEAA
| IBCCBF2F5A49A76D461A7479DA2813EA7 | IABDBB85ACD3277D447B4FD8665EA150B | IEB1DC53BA14A2028F346A4C10651DA08 ; assign
IB624795CEFFC2094E111CAD5578DAE1C = I95628D4658FCAB1EADD1EBA1F6294ED6 | I2A46DB8D4D31FAC435A47D582BA0E704 | IB55475954FE95F83F22B1C2FB76FAEC7
| I38BDB4EBCC779338E7AF863601C4853E | I270710745C28824E285C2E05FB618D27 | IFFE90484B4E519D0DD55AFC0D9379B2A | IB77F87CED77CEC2F6256375F35443CD0
| I7616B3B0828958A3CA36203B840CF4D6 ; assign IB56580C539321C40E6B44EB394A9EECF = I841AB9A2043753D035FC3A85DEFAF1D2
| IF6683BD4A4C0331D12A89BC5CD3FDAA2 | I31980ABC07D19BA89784085C7754DE42 | ICD34F2C7357A369358E7CFBC3D425106 | I765A5C6CB6D2AE7496EF2BE962529E09
| I6FDDB4608592CC601F82E29CF03F58E2 | IAF3303768435E5C76A60A5987AF1CD0A | I246B1D75EEA1239D65C20304AF791CB4 ; assign
I400149787F2546E3D0331041FB8123FC = {IBCEA86C0BDF1E124E6697E40D620DD0A , I2130A737A8CF0DAA0688CD61C692C53A , IE6E0B2D716FF39D4E07D15E9EAAB04FC ,
I9C559D18449178998B7475813A7D0CBB , I081CFEF0428EFE96BD06A8F2EE9DC2CD , IE1F9397E899B4E938A0D54FC51445C13 , I40DCE993F9A1E526661825B1281A7DCB ,
I711EA37894AB982C997C1497E71677B4 }; assign I97E631353C4C7709CF07D5FC5800DDBC = I42DFCF8044FC66463EFBDCD6F2C69AEE
| I9A3A1B70A9C668CF11493348B519FF4B | IDE0F2D42601304C0E0CCD60778B3938F | ID34187ADCB71E296DE727A7573E76A15 | I7B62DE436B5B4C0A20CC4FE1E5D6F91D
| IA2F68AF483F09457F392B22939441F47 | I009BA1F74DBCC8E4177F1254D60DCAE9 | I11D20DB2F186022215040429BE705A72 ; assign
I56519DD369C66F1A0EA1EE3D2398E0EF = {I8824AFA21C1B61513D8DE94591B948FB , IE67F175E6F2CC66DDCAD62CCD21F3551 , IE0683883BF201CF74ADDEE61816AAD96 ,
I82635882370B55739EA7454635CE3A41 , IA3A543EBA3F35D293D9F9A372241FFB7 , I3ABE7E8A0A3ADCF18D9C06A84D938210 , I5B92AFCE2F6F881BA10FA726B18BB692 ,
I6FE2694F3F3B5838177CEF5992A016F2 , I6AF9911F8AAC2F653011D5D8ACE5F433 }; assign IC0667A37FE3E5F8D3579C6AEF86F5C24
= {IB5292E1DAB3B0E7E62E43F792E80D8F1 , {8{1'b0}}}; assign IED75BA58ED5F09B80AEBB5C4531DD96E = I6DFBACFF2E5A466B93A00001848429F7
| I49850943EA73C8BE46401A2FC9B67D74 | I386D96EE2FCEC8374B24F3017B94BD4D | I98308209671212A3C88A9644B503FA02 | I88DEF602C28E2AE7FCFC75761E9DF8F6
| I0D8A716B0016AFE64E7F7977A80A253A | IFFB9EED620356BDFB94697DB3606174F | I3E4C4B769B824746306BEC19D75E1A23 | I1179A173C6F4C43BA9C3B71086E48486 ;
assign I86E103F0E5684240BF4D6AD4E9635C7A = I7CA41EFBA3D0548B989711570EA40B95 | I14F6DF0BCAC12F6EBAD7145BDD4B2D26
| I11E1C086CA3C13B481A5977B8AD8694F | IB4C822D6BFAE40F12254437B18142B8A | I6434FE6B1DB9B4DCDB82F1E568D8A5AD | IAEFBAA4728FB6854C056C8E4C0691B3D
| I2C072E656BFCADF4877B42244D6D2307 | IA2B524351B6A8AB3A2FA7E1B456ABE67 | IC99E8E0D5BAC180B4FAC3C67D1618142 ; assign
I6618736D0C53F4C6D20F8C252BF264AD = IC30C68A9857DD63CE5A51E5943CEB3AF | IB85FB30E34AF0B105FD21BBBB73605EA | I5C58E3085FDB240D9A5DD64A9CD3A30B
| I30157CAB406F288B630EF42C05ACC134 | IF76FEAB2FA7E91BC33928D6B232B6040 | I1DC328E1B03775141AFCFBB60C78CDC0 | IB96A9322FAF5941DF70737CA69F152A3
| I037B294714AE918C1D513F83470C0190 | I1C08DD68F49BF5FFE04D852950D9A932 ;  generate begin if (IA54DA90446D375855AF33292D2570A3C )
for (I24501E622BFA6932719D2F78F75F6270 = 0; I24501E622BFA6932719D2F78F75F6270 < 32; I24501E622BFA6932719D2F78F75F6270
= I24501E622BFA6932719D2F78F75F6270 + 1) if (I24501E622BFA6932719D2F78F75F6270 < IA54DA90446D375855AF33292D2570A3C )
assign I97B15B5DA5A0868F11CDF3929B25044E [I24501E622BFA6932719D2F78F75F6270 ] = I1C0271AD5E8E9E9164909E468AD0B212 [I24501E622BFA6932719D2F78F75F6270 ];
else assign I97B15B5DA5A0868F11CDF3929B25044E [I24501E622BFA6932719D2F78F75F6270 ] = 1'b0; else assign I97B15B5DA5A0868F11CDF3929B25044E
= 32'b0; end endgenerate generate begin if (IE50492CEE03959C13AD5E521CC7F2FEF && (I97F18A3381F2546EB21E07DF7628912F
> 0)) for (I24501E622BFA6932719D2F78F75F6270 = 0; I24501E622BFA6932719D2F78F75F6270 < 32; I24501E622BFA6932719D2F78F75F6270
= I24501E622BFA6932719D2F78F75F6270 + 1) if (I24501E622BFA6932719D2F78F75F6270 < I97F18A3381F2546EB21E07DF7628912F )
assign I16A1A5B65742A57E7143E981BF286F99 [I24501E622BFA6932719D2F78F75F6270 ] = I1C0271AD5E8E9E9164909E468AD0B212 [IA54DA90446D375855AF33292D2570A3C
+ I24501E622BFA6932719D2F78F75F6270 ]; else assign I16A1A5B65742A57E7143E981BF286F99 [I24501E622BFA6932719D2F78F75F6270 ]
= 1'b0; else assign I16A1A5B65742A57E7143E981BF286F99 = 32'b0; end endgenerate generate begin if (I0B3C14F69FAC563649E26679A3D8B1CD
&& (I0069A39965C0330678D64B612F60F78D > 0)) for (I24501E622BFA6932719D2F78F75F6270 = 0; I24501E622BFA6932719D2F78F75F6270
< 32; I24501E622BFA6932719D2F78F75F6270 = I24501E622BFA6932719D2F78F75F6270 + 1) if (I24501E622BFA6932719D2F78F75F6270
< I0069A39965C0330678D64B612F60F78D ) assign IB4CA57E47B085EE5925036D5223A4598 [I24501E622BFA6932719D2F78F75F6270 ]
= I1C0271AD5E8E9E9164909E468AD0B212 [IA54DA90446D375855AF33292D2570A3C + I97F18A3381F2546EB21E07DF7628912F + I24501E622BFA6932719D2F78F75F6270 ];
else assign IB4CA57E47B085EE5925036D5223A4598 [I24501E622BFA6932719D2F78F75F6270 ] = 1'b0; else assign IB4CA57E47B085EE5925036D5223A4598
= 32'b0; end endgenerate generate begin if (IFA272F301A5935EE15CB134524665363 && (IC69BEB80DB094A65F3DFB0265F8616DE
> 0)) for (I24501E622BFA6932719D2F78F75F6270 = 0; I24501E622BFA6932719D2F78F75F6270 < 32; I24501E622BFA6932719D2F78F75F6270
= I24501E622BFA6932719D2F78F75F6270 + 1) if (I24501E622BFA6932719D2F78F75F6270 < IC69BEB80DB094A65F3DFB0265F8616DE )
assign I2F92739468FA7128C93936C8511AA228 [I24501E622BFA6932719D2F78F75F6270 ] = I1C0271AD5E8E9E9164909E468AD0B212 [IA54DA90446D375855AF33292D2570A3C
+ I97F18A3381F2546EB21E07DF7628912F + I0069A39965C0330678D64B612F60F78D + I24501E622BFA6932719D2F78F75F6270 ]; else
assign I2F92739468FA7128C93936C8511AA228 [I24501E622BFA6932719D2F78F75F6270 ] = 1'b0; else assign I2F92739468FA7128C93936C8511AA228
= 32'b0; end endgenerate generate begin if (IE690B7723F136DA02896C0728DDADB49 && (I4046611EA3EEF60ACE26738C818FDBA2
> 0)) for (I24501E622BFA6932719D2F78F75F6270 = 0; I24501E622BFA6932719D2F78F75F6270 < 32; I24501E622BFA6932719D2F78F75F6270
= I24501E622BFA6932719D2F78F75F6270 + 1) if (I24501E622BFA6932719D2F78F75F6270 < I4046611EA3EEF60ACE26738C818FDBA2 )
assign I25DCCEF37BE2FCC042C00B81ABCA449F [I24501E622BFA6932719D2F78F75F6270 ] = I1C0271AD5E8E9E9164909E468AD0B212 [IA54DA90446D375855AF33292D2570A3C
+ I97F18A3381F2546EB21E07DF7628912F + I0069A39965C0330678D64B612F60F78D + IC69BEB80DB094A65F3DFB0265F8616DE + I24501E622BFA6932719D2F78F75F6270 ];
else assign I25DCCEF37BE2FCC042C00B81ABCA449F [I24501E622BFA6932719D2F78F75F6270 ] = 1'b0; else assign I25DCCEF37BE2FCC042C00B81ABCA449F
= 32'b0; end endgenerate generate begin if (I55BE27080C370AF723A4FE096014E875 && (IAE03DAE231BA40E8DD1C02D38068EF8A
> 0)) for (I24501E622BFA6932719D2F78F75F6270 = 0; I24501E622BFA6932719D2F78F75F6270 < 32; I24501E622BFA6932719D2F78F75F6270
= I24501E622BFA6932719D2F78F75F6270 + 1) if (I24501E622BFA6932719D2F78F75F6270 < IAE03DAE231BA40E8DD1C02D38068EF8A )
assign I19381BD04F07A020B45A7EFE952EBD90 [I24501E622BFA6932719D2F78F75F6270 ] = I1C0271AD5E8E9E9164909E468AD0B212 [IA54DA90446D375855AF33292D2570A3C
+ I97F18A3381F2546EB21E07DF7628912F + I0069A39965C0330678D64B612F60F78D + IC69BEB80DB094A65F3DFB0265F8616DE + I4046611EA3EEF60ACE26738C818FDBA2
+ I24501E622BFA6932719D2F78F75F6270 ]; else assign I19381BD04F07A020B45A7EFE952EBD90 [I24501E622BFA6932719D2F78F75F6270 ]
= 1'b0; else assign I19381BD04F07A020B45A7EFE952EBD90 = 32'b0; end endgenerate generate begin if (IB2560D175E4507798B84D6E659FD6373
&& (I7568F6D9A53738CCE095CE231BAB3F85 > 0)) for (I24501E622BFA6932719D2F78F75F6270 = 0; I24501E622BFA6932719D2F78F75F6270
< 32; I24501E622BFA6932719D2F78F75F6270 = I24501E622BFA6932719D2F78F75F6270 + 1) if (I24501E622BFA6932719D2F78F75F6270
< I7568F6D9A53738CCE095CE231BAB3F85 ) assign ID54A2FD9EE0AEAC4E7AC2A4D30D28B9B [I24501E622BFA6932719D2F78F75F6270 ]
= I1C0271AD5E8E9E9164909E468AD0B212 [IA54DA90446D375855AF33292D2570A3C + I97F18A3381F2546EB21E07DF7628912F + I0069A39965C0330678D64B612F60F78D
+ IC69BEB80DB094A65F3DFB0265F8616DE + I4046611EA3EEF60ACE26738C818FDBA2 + IAE03DAE231BA40E8DD1C02D38068EF8A + I24501E622BFA6932719D2F78F75F6270 ];
else assign ID54A2FD9EE0AEAC4E7AC2A4D30D28B9B [I24501E622BFA6932719D2F78F75F6270 ] = 1'b0; else assign ID54A2FD9EE0AEAC4E7AC2A4D30D28B9B
= 32'b0; end endgenerate generate begin if (I25B649490B20A1FEC9A1AA60AB0C6D5E && (IEB4CAA0AE4F26FAC1DAA6B9884179DEA
> 0)) for (I24501E622BFA6932719D2F78F75F6270 = 0; I24501E622BFA6932719D2F78F75F6270 < 32; I24501E622BFA6932719D2F78F75F6270
= I24501E622BFA6932719D2F78F75F6270 + 1) if (I24501E622BFA6932719D2F78F75F6270 < IEB4CAA0AE4F26FAC1DAA6B9884179DEA )
assign IA5469486BB0530B9AA1B819A3C7A9583 [I24501E622BFA6932719D2F78F75F6270 ] = I1C0271AD5E8E9E9164909E468AD0B212 [IA54DA90446D375855AF33292D2570A3C
+ I97F18A3381F2546EB21E07DF7628912F + I0069A39965C0330678D64B612F60F78D + IC69BEB80DB094A65F3DFB0265F8616DE + I4046611EA3EEF60ACE26738C818FDBA2
+ IAE03DAE231BA40E8DD1C02D38068EF8A + I7568F6D9A53738CCE095CE231BAB3F85 + I24501E622BFA6932719D2F78F75F6270 ]; else
assign IA5469486BB0530B9AA1B819A3C7A9583 [I24501E622BFA6932719D2F78F75F6270 ] = 1'b0; else assign IA5469486BB0530B9AA1B819A3C7A9583
= 32'b0; end endgenerate  I2296FC491415818D18357D6C2D700C14 # ( .IFC1FF746397E6A576E9FEB281890A248 (I857673E5DE2CF777499EE369473CBCCC ),
.IAF1DF965ED0D670C125D16FDF91B875B (IA874AED52F9C16F13B580898DA0E85AC ), .IB7B379BA36F36F0638F4F33C7598CC85 (I45E74A319CD545DA84EE876844F12DF8 ),
.ID9DCCEB6B5B42C479CB9D2B3C992035D (I212658651766EFCF73257AF1E3121AF8 ), .I251C6E5612F7B344EC3156CB9A93BE5B (I2610FF174BEEE098C8D9C9374191F122 ),
.ID7A688D3DA9A2C539FE87FC8998248CB (IA8729443C3DAFAFDD37A6BED4B24F26C ), .I96DBC3D130FB2B57DFB76E3E87DF89D2 (I08EC85B0527EBF111FDA96E4BD71B6BF ),
.I87B53E44EDBDCDA1796FB105323D3B17 (I6C75B7796A1597A63620710B69C04958 ), .IF9554E0938E353BDC05ABE0C628E3BE9 (I86AD8EB6B8FA8A1AA6EA64DE4357E4EA ),
.I37C708634F442A3B0568DA0BB576511F (I5C0FF6EA47D5544D48B9200C35F2015D ), .I7B125DA60401B7C86EB027E9E9262847 (IED6EFA8FE915B71B8E198535343CFBFB ),
.I8BEE88809FA5712893BC59FF0E17ADB2 (I98F26EACDFB5625667BCAFBDB2867748 ), .I7DF5A90920A562D09AA22D2DFA657124 (I3CAEAE4A6B7BA30F88F0945373893582 ),
.I0243B4A4E84E0712929C806F438E6AA9 (ICC1064DA289312A92936196EA26F0023 ), .I7050B96C0C45A812BBFC45C2A30F272C (I78F9B7090517BBEEBC1543199FBA4D34 ),
.IB7C70D5D7B0DDF146F4D402BEE6F6FA6 (I731C578B2B8A6173399D3CABA7E98889 ), .I1CBD8B214B4765FBC7FA828F0C62BC94 (IE18DEDE16538C154B2EFCB2652C25FD5 ),
.I677BE3663880CBE6E5AE2C431F3FDD4D (IB6EB169241E23C32C11DDDC27322BCE6 ), .I1CF1EE9FA60C0CDB15DD404CC8A269E5 (I83476C8D11033DBF952882C55FC0E55B ),
.I34F020684BFF4B1EAA406E693751B71D (I156838D82D20DC7C269685B24CB4A8B0 ), .IFB94B817F0BC84EC0734110F6EDE475A (I86134D1B828E3E59B9C4B66EC0920D98 ),
.I512A575E055CF9235066DBE4051242CB (IC2EB58967FBD1CD5C54491738F4BAD86 ), .I391BF6A9C9F2ABEEA227F0E1F3F50A4F (IBBBF11BAEEC8458B08DFB6E2D9D1C850 ),
.IF0D7F78B99E50997A728E3731A197225 (IA54DA90446D375855AF33292D2570A3C ), .I9606837003EFA36A64A97C352D3D89A3 (IAD54DD4DF3ABBB4563A2B75498325CD7 ),
.I4C1994114E1C49B9376320858F4E71F9 (I02756A8C58D5B37B7049B7F6FA2073B7 ), .I2CB8399B2A61CDA9DB269D3567018E65 (I1066D287D755AADD24EE379E400F8DA8 ),
.I46C5269B9FB24EF04CE2CC341C288EC7 (I46C5269B9FB24EF04CE2CC341C288EC7 ), .I3C9AD458B89B2FAABD743BF4E13BF421 (I3C9AD458B89B2FAABD743BF4E13BF421 ),
.I73ABD5619A9FB885445AC1E288EAF7F8 (0), .IBDE0431C8F903800F409661F4F56FD80 (IB26EBF559CA483EACBAD1BCA4C580AF2 )
) IA2EA3BC627C5D679C3AE5BCC26B64F6D ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .ICB680FEAB46B6D635CD9DD6BB49A6A20 (IEE7B9D1B054F5CACBC10351FC32D7BFA ), .I8FF768DAF4C56D1B2D217B2C02B6D4EC
(IFE8155182FD754C22D6F7FDA1F1C1174 ), .I9E5E6E86745F53F982BC3862031A206B (ICFA3AEC9D2E8697060447D8D8EB18A80 ), .I3AD72E1D6C16169DB8A27F1681293009
(I81D61D198832883CFD88EB5DEB88A32B ), .I0DE44F162EF92573C5DE1249527F6E9D (I1F5A786F105B576AC15A6F25EBFB89B8 ), .I2E9CC9AFC2E4742F852CB037CFC7E0A1
(IB9B532CA44CE4054811AB748EDD0922D ), .I8B1798242C3B0E655181D0D365813614 (I8B1798242C3B0E655181D0D365813614 ), .IE145222FDBDC80109E12FA72D3D3C655
(IE145222FDBDC80109E12FA72D3D3C655 ), .ID43AC1009727D128F1C5DFE4640CA5AB (ID43AC1009727D128F1C5DFE4640CA5AB ), .IB610431939CB8180EAC2403672BAF58D
(IB610431939CB8180EAC2403672BAF58D ), .I3C7A9FA839F554D8898020C4831479E2 (IC7DB18773990D347CEF55E672D6B2C05 ), .I74A0936EE8FD1443A2C6745A4F3F6B5E
(I39A06B46F4E1C11EE4BFB781E3B4F32A ), .I369BA2FFB5D41DF25F9BC3AB126D6607 (I369BA2FFB5D41DF25F9BC3AB126D6607 ), .I1C0271AD5E8E9E9164909E468AD0B212
(I97B15B5DA5A0868F11CDF3929B25044E ), .I6EC1BE4B18EC6AA3D88A5D45B614565E (I6EC1BE4B18EC6AA3D88A5D45B614565E [0]),
.I56148DDDF284443347FFCF4F9C3BE61A (I81BF37FCB51B492DCA857F28ABD8D76E [0]), .I24C403550AE065D7D1B7266142886226 (I24C403550AE065D7D1B7266142886226 ),
.I438B8BD876741F9B46EB770E92F808B7 (I438B8BD876741F9B46EB770E92F808B7 [11:0]), .I5FE75BE614D4F52DB327549B36203350
(I74CF4D6FE5B30BB30E40AFCA2A08A220 [0]), .I3D6C771D05CA1A769E61302C086494B8 (I3D6C771D05CA1A769E61302C086494B8 ),
.I357B3043EDACE3EBECE8F54D79B9F90A (I357B3043EDACE3EBECE8F54D79B9F90A ), .I0AAD559CF33A5CBA597990658774FEB3 (I0AAD559CF33A5CBA597990658774FEB3 ),
.I923204A95D8CBB206587CF32BEDCF4EF (I923204A95D8CBB206587CF32BEDCF4EF ), .ICF9D8FD31DFC7D20DAF939C6D75F1518 (ICF9D8FD31DFC7D20DAF939C6D75F1518 [0]),
.IDF550B17734BF16B7E410B19BB31E276 (I5917F25EB5F020E0FEEB03EB956B3110 ), .I8ED9B9C1D9F58C5D06A9443AD901E8C6 (I9818F0A46507B01B5AAD29ECB3D36F81 ),
.IA976D63BEECA80DCE31365CF56EC0248 (I0EB153824311AB3255F80A6B20F59828 ), .I5E3CE5AF5C34D232BFB139B63D9912B4 (I6A77961ADE4327F78C7D008C5DA7D184 ),
.IBEF3E5F9395E2C7822AE03D6461DEBBB (I8C1666B519246534E1C4722652FD1823 ), .I7E6CFD6A7DCAB9CD2188D044C7D716A6 (I95628D4658FCAB1EADD1EBA1F6294ED6 ),
.I3A34691662384260F0524DD7F650E75A (I841AB9A2043753D035FC3A85DEFAF1D2 ), .IC2F58AB5028C1D2C53C6EF47A4975D0A (I711EA37894AB982C997C1497E71677B4 ),
.I112E0A79129A8BC6DD4C13647C31F8A0 (I42DFCF8044FC66463EFBDCD6F2C69AEE ), .IE4B6DD43E04940631EF58BA04EA58997 (IACF97B89AE62537A26788BDFCE846ED1 [0]),
.I3A095084CDFDFA56A0E67616A78D3B25 (I01D4C6B20466D26621C6DA5816817455 [0]), .I81CD7F184DF8D58A1F2324E975A6816C (I46A701488EBE724B47736C3C7A47A876 [0]),
.I83C4A4200EB2B3F6766D338284ECAAAF (IFE63F76C2A46B87271596BE8D0FFD21A [0]), .I42A419EB6EB8D11234AC3B2BCA0AE593 (I999118EB4E0839ECF8CF049C93027B49 ),
.IA41AC3CC6BC050DDC172724AB311315B (I6080D873E932E26F13608A1D73FAE7C0 ), .I31CF69FF368B36B4D6612DF16B3ABC6B (I21EE6CA5EBC86B66AC5EE8AF763FB838 [0]),
.IFE4A8CBA73734C6F0F0A078027E053D4 (I1179A173C6F4C43BA9C3B71086E48486 ), .ID7A2A8B1E9D92B60194D5FAFAAB15208 (IC99E8E0D5BAC180B4FAC3C67D1618142 ),
.IF274FAF97F5BACD693913BB418717A9D (I1C08DD68F49BF5FFE04D852950D9A932 ), .ID95C13E7EE1CFE6A8743FF9E62C25873 (I6AF9911F8AAC2F653011D5D8ACE5F433 ),
.IC58E411F24D810EF60A7B8638ABCC0BB (I7D2B5C97BC25D475F870C1BE7E21B697 ), .I89CFFA73C7546481B72B0FB06D799AEE (IF082298B35C4A83318C3597AC50DA20E ),
.I270ED686C2EF2C1C8B5B55EC4A5AAE84 (I762EB11F447E9FE5C306D10B1D44F3D1 ), .ID5CCD4858CB5CC1B2EDEC682C7DE5AAD (I7ED71D3164ABC636AC5046B7E263FD03 ),
.I7D901091F9E0741061C75B54467D48A0 (I6795B29551221467FFA6B7172DDA857D ) );  generate if (IE50492CEE03959C13AD5E521CC7F2FEF )
I2296FC491415818D18357D6C2D700C14 # ( .IFC1FF746397E6A576E9FEB281890A248 (IE8C1215A45516D3178A8A93152E05EE2 ), .IAF1DF965ED0D670C125D16FDF91B875B
(I6A67F4FE467D33BBE90E5158D72171A4 ), .IB7B379BA36F36F0638F4F33C7598CC85 (I8F998DCDBE9627EA583F7BB408EC780D ), .ID9DCCEB6B5B42C479CB9D2B3C992035D
(I8695C513BA5D9DA307CC481D6AFFB133 ), .I251C6E5612F7B344EC3156CB9A93BE5B (IEE21CD471C5E4E6CE83A164513BC7722 ), .ID7A688D3DA9A2C539FE87FC8998248CB
(I56DA37D670BDECB81356B81560DC8649 ), .I96DBC3D130FB2B57DFB76E3E87DF89D2 (IB36C0E6BB9CF8D4E4A2F31086369A6EC ), .I87B53E44EDBDCDA1796FB105323D3B17
(I6C4BB963A9FEECAA07E250007DE29E69 ), .IF9554E0938E353BDC05ABE0C628E3BE9 (I7725F462040C54BFDFC296100F95D5D0 ), .I37C708634F442A3B0568DA0BB576511F
(IC022347DC0BBA44450EA061654CE4130 ), .I7B125DA60401B7C86EB027E9E9262847 (I8DFF460C39C720D8E01DF9AD54E62457 ), .I8BEE88809FA5712893BC59FF0E17ADB2
(I128970AF889EC52F4195C246A49524BA ), .I7DF5A90920A562D09AA22D2DFA657124 (I61E4D6D4FFCCB1C283902514C76CD3AA ), .I0243B4A4E84E0712929C806F438E6AA9
(ID0832173F4D69F0B96DB00FA9805F75F ), .I7050B96C0C45A812BBFC45C2A30F272C (I171E938E7CDE23987F02EB923184A5C3 ), .IB7C70D5D7B0DDF146F4D402BEE6F6FA6
(I5A509B803B47567D6FA4F4CB4C6AA95D ), .I1CBD8B214B4765FBC7FA828F0C62BC94 (I2C1FDD71B618A0C398964466A5958BF0 ), .I677BE3663880CBE6E5AE2C431F3FDD4D
(ICE7C691E1DC04B92371B76DCE234C732 ), .I1CF1EE9FA60C0CDB15DD404CC8A269E5 (IA9D9F2D7EEC92A228D6CC71EE9A86E0E ), .I34F020684BFF4B1EAA406E693751B71D
(I7356A0718B40AEF099CE99273A8CBC19 ), .IFB94B817F0BC84EC0734110F6EDE475A (I4521B8E3C71C6E5D7639756B81D56C58 ), .I512A575E055CF9235066DBE4051242CB
(IB52E64F4A5E8239ED2BF949AC0702ACE ), .I391BF6A9C9F2ABEEA227F0E1F3F50A4F (IA5A53C930B674A8F9761966972CFB6F6 ), .IF0D7F78B99E50997A728E3731A197225
(I97F18A3381F2546EB21E07DF7628912F ), .I9606837003EFA36A64A97C352D3D89A3 (I2FCDB5B825200EDE4D7757A0621663E0 ), .I4C1994114E1C49B9376320858F4E71F9
(IC745524098FFC5FBA778DA59D2444D9B ), .I2CB8399B2A61CDA9DB269D3567018E65 (I7507C2B666C444A66EDA2CFDB6DCEEB9 ), .I46C5269B9FB24EF04CE2CC341C288EC7
(I46C5269B9FB24EF04CE2CC341C288EC7 ), .I3C9AD458B89B2FAABD743BF4E13BF421 (I3C9AD458B89B2FAABD743BF4E13BF421 ), .I73ABD5619A9FB885445AC1E288EAF7F8
(1), .IBDE0431C8F903800F409661F4F56FD80 (IB26EBF559CA483EACBAD1BCA4C580AF2 ) ) I6783E3B3DCEAE9D0ED0773BD1B72AC00
( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ),
.ICB680FEAB46B6D635CD9DD6BB49A6A20 (I7FE73B332A2A7E273F8EC82CC2A0A9D1 ), .I8FF768DAF4C56D1B2D217B2C02B6D4EC (I8C784B1A25E6B5F5402709647F921D20 ),
.I9E5E6E86745F53F982BC3862031A206B (IAFB7D4809B407BA0A70ABF120DF37844 ), .I3AD72E1D6C16169DB8A27F1681293009 (IA69AD6BF563BE83DB737C644B2992470 ),
.I0DE44F162EF92573C5DE1249527F6E9D (IBBC01C0CF0EE486327FBEB391C90772B ), .I2E9CC9AFC2E4742F852CB037CFC7E0A1 (I147607D1A744B7E8E0F3050C499F3A23 ),
.I8B1798242C3B0E655181D0D365813614 (I8B1798242C3B0E655181D0D365813614 ), .IE145222FDBDC80109E12FA72D3D3C655 (IE145222FDBDC80109E12FA72D3D3C655 ),
.ID43AC1009727D128F1C5DFE4640CA5AB (ID43AC1009727D128F1C5DFE4640CA5AB ), .IB610431939CB8180EAC2403672BAF58D (IB610431939CB8180EAC2403672BAF58D ),
.I3C7A9FA839F554D8898020C4831479E2 (IC7DB18773990D347CEF55E672D6B2C05 ), .I74A0936EE8FD1443A2C6745A4F3F6B5E (I39A06B46F4E1C11EE4BFB781E3B4F32A ),
.I369BA2FFB5D41DF25F9BC3AB126D6607 (I369BA2FFB5D41DF25F9BC3AB126D6607 ), .I1C0271AD5E8E9E9164909E468AD0B212 (I16A1A5B65742A57E7143E981BF286F99 ),
.I6EC1BE4B18EC6AA3D88A5D45B614565E (I6EC1BE4B18EC6AA3D88A5D45B614565E [1]), .I56148DDDF284443347FFCF4F9C3BE61A (I81BF37FCB51B492DCA857F28ABD8D76E [1]),
.I24C403550AE065D7D1B7266142886226 (I24C403550AE065D7D1B7266142886226 ), .I438B8BD876741F9B46EB770E92F808B7 (I438B8BD876741F9B46EB770E92F808B7 [11:0]),
.I5FE75BE614D4F52DB327549B36203350 (I74CF4D6FE5B30BB30E40AFCA2A08A220 [1]), .I3D6C771D05CA1A769E61302C086494B8 (I3D6C771D05CA1A769E61302C086494B8 ),
.I357B3043EDACE3EBECE8F54D79B9F90A (I357B3043EDACE3EBECE8F54D79B9F90A ), .I0AAD559CF33A5CBA597990658774FEB3 (I0AAD559CF33A5CBA597990658774FEB3 ),
.I923204A95D8CBB206587CF32BEDCF4EF (I923204A95D8CBB206587CF32BEDCF4EF ), .ICF9D8FD31DFC7D20DAF939C6D75F1518 (ICF9D8FD31DFC7D20DAF939C6D75F1518 [1]),
.IDF550B17734BF16B7E410B19BB31E276 (I25D510B1A7EEBD7D688C48A4050B0A28 ), .I8ED9B9C1D9F58C5D06A9443AD901E8C6 (I85BF4AD7C60BEA5045D19571D851C992 ),
.IA976D63BEECA80DCE31365CF56EC0248 (IBF1BA20BCDFE79989AD3C8104A1024A4 ), .I5E3CE5AF5C34D232BFB139B63D9912B4 (I4B2CDC61C9F80778CDBA134570DB93A1 ),
.IBEF3E5F9395E2C7822AE03D6461DEBBB (IB3122CB8FBD2C123E9D9BD0599AE41D0 ), .I7E6CFD6A7DCAB9CD2188D044C7D716A6 (I2A46DB8D4D31FAC435A47D582BA0E704 ),
.I3A34691662384260F0524DD7F650E75A (IF6683BD4A4C0331D12A89BC5CD3FDAA2 ), .IC2F58AB5028C1D2C53C6EF47A4975D0A (I40DCE993F9A1E526661825B1281A7DCB ),
.I112E0A79129A8BC6DD4C13647C31F8A0 (I9A3A1B70A9C668CF11493348B519FF4B ), .IE4B6DD43E04940631EF58BA04EA58997 (IACF97B89AE62537A26788BDFCE846ED1 [1]),
.I3A095084CDFDFA56A0E67616A78D3B25 (I01D4C6B20466D26621C6DA5816817455 [1]), .I81CD7F184DF8D58A1F2324E975A6816C (I46A701488EBE724B47736C3C7A47A876 [1]),
.I83C4A4200EB2B3F6766D338284ECAAAF (IFE63F76C2A46B87271596BE8D0FFD21A [1]), .I42A419EB6EB8D11234AC3B2BCA0AE593 (I09A93891DA1B4315581C9B6775306EC6 ),
.IA41AC3CC6BC050DDC172724AB311315B (IA60C7697AAB3A707DC265C02AA59526E ), .I31CF69FF368B36B4D6612DF16B3ABC6B (I21EE6CA5EBC86B66AC5EE8AF763FB838 [1]),
.IFE4A8CBA73734C6F0F0A078027E053D4 (I3E4C4B769B824746306BEC19D75E1A23 ), .ID7A2A8B1E9D92B60194D5FAFAAB15208 (IA2B524351B6A8AB3A2FA7E1B456ABE67 ),
.IF274FAF97F5BACD693913BB418717A9D (I037B294714AE918C1D513F83470C0190 ), .ID95C13E7EE1CFE6A8743FF9E62C25873 (I6FE2694F3F3B5838177CEF5992A016F2 ),
.IC58E411F24D810EF60A7B8638ABCC0BB (I976ABC47C39290CF3E29B8773D338ECE ), .I89CFFA73C7546481B72B0FB06D799AEE (I42864A73C6A7A061BF0E25880AF8AE9C ),
.I270ED686C2EF2C1C8B5B55EC4A5AAE84 (I24FB1AC5C4A1C96F7DF559EABAD558C5 ), .ID5CCD4858CB5CC1B2EDEC682C7DE5AAD (ICA544D75FD0BAE421ECEFDBC4207F6C1 ),
.I7D901091F9E0741061C75B54467D48A0 (IEC017B3AB9F16AE871D5253A5257D941 ) ); else begin assign ICF9D8FD31DFC7D20DAF939C6D75F1518 [1]
= 1'b0; assign IACF97B89AE62537A26788BDFCE846ED1 [1] = 1'b0; assign I01D4C6B20466D26621C6DA5816817455 [1] = 1'b0;
assign I46A701488EBE724B47736C3C7A47A876 [1] = 1'b0; assign IFE63F76C2A46B87271596BE8D0FFD21A [1] = 1'b0; assign
I21EE6CA5EBC86B66AC5EE8AF763FB838 [1] = 1'b0; assign I25D510B1A7EEBD7D688C48A4050B0A28 = 1'b0; assign I85BF4AD7C60BEA5045D19571D851C992
= 1'b0; assign IBF1BA20BCDFE79989AD3C8104A1024A4 = 1'b0; assign I4B2CDC61C9F80778CDBA134570DB93A1 = 1'b0; assign
IB3122CB8FBD2C123E9D9BD0599AE41D0 = 1'b0; assign I2A46DB8D4D31FAC435A47D582BA0E704 = 1'b0; assign IF6683BD4A4C0331D12A89BC5CD3FDAA2
= 1'b0; assign I40DCE993F9A1E526661825B1281A7DCB = 1'b0; assign I9A3A1B70A9C668CF11493348B519FF4B = 3'b0; assign
I09A93891DA1B4315581C9B6775306EC6 = 3'b0; assign IA60C7697AAB3A707DC265C02AA59526E = 3'b0; assign I3E4C4B769B824746306BEC19D75E1A23
= 32'b0; assign IA2B524351B6A8AB3A2FA7E1B456ABE67 = 1'b0; assign I037B294714AE918C1D513F83470C0190 = 1'b0; assign
I6FE2694F3F3B5838177CEF5992A016F2 = 1'b0; assign I976ABC47C39290CF3E29B8773D338ECE = 11'b0; assign I42864A73C6A7A061BF0E25880AF8AE9C
= 1'b0; assign I24FB1AC5C4A1C96F7DF559EABAD558C5 = 1'b0; assign ICA544D75FD0BAE421ECEFDBC4207F6C1 = 1'b0; assign
IEC017B3AB9F16AE871D5253A5257D941 = 32'b0; end endgenerate  generate if (I0B3C14F69FAC563649E26679A3D8B1CD ) I2296FC491415818D18357D6C2D700C14
# ( .IFC1FF746397E6A576E9FEB281890A248 (I1A39FC80F18CFB225DD25F1158A43FEB ), .IAF1DF965ED0D670C125D16FDF91B875B
(IFA1CC1A50C8D64B9481E806D15AF3CA5 ), .IB7B379BA36F36F0638F4F33C7598CC85 (IF089B8BB6C2663DE1CA53AB4AB67231B ), .ID9DCCEB6B5B42C479CB9D2B3C992035D
(I348F387B0CC3540AF0215535F676D5A2 ), .I251C6E5612F7B344EC3156CB9A93BE5B (I3AB6DCBD252A38D5954C33DB9CFA020B ), .ID7A688D3DA9A2C539FE87FC8998248CB
(IFE55C92252D5A4FCF3878CC98FCAD612 ), .I96DBC3D130FB2B57DFB76E3E87DF89D2 (IC2181A40E4750EEA118AA81ABB4E415B ), .I87B53E44EDBDCDA1796FB105323D3B17
(I813CE6D8049DC9123C58691D1DA81B59 ), .IF9554E0938E353BDC05ABE0C628E3BE9 (I50243AFBCB64F92A3F6EEC157034F4FC ), .I37C708634F442A3B0568DA0BB576511F
(I38E6C6DF2535A2049746702855108B5A ), .I7B125DA60401B7C86EB027E9E9262847 (I0FFEAFBF23F15260885D040F12B66960 ), .I8BEE88809FA5712893BC59FF0E17ADB2
(I31E80F0EE05B52A92941F617BDCEF890 ), .I7DF5A90920A562D09AA22D2DFA657124 (I509611AF740C942BA82FB9ECE7BA4E67 ), .I0243B4A4E84E0712929C806F438E6AA9
(I586C95E6CCC79680B179527AE8977C4E ), .I7050B96C0C45A812BBFC45C2A30F272C (I39D41D0CFF63339D485BDBCDBC3A8729 ), .IB7C70D5D7B0DDF146F4D402BEE6F6FA6
(IF833CBC3D7A215E6C5635F3F07A09365 ), .I1CBD8B214B4765FBC7FA828F0C62BC94 (IE106099B16008BAE163236DC5CF4EAFE ), .I677BE3663880CBE6E5AE2C431F3FDD4D
(IC4C3CD51A29DC2F222334D23407BB4E7 ), .I1CF1EE9FA60C0CDB15DD404CC8A269E5 (I7C988FF99F8B28AB1CE2299774306236 ), .I34F020684BFF4B1EAA406E693751B71D
(I4FF1FE282379DCB83A2AF4F7A12AF6CA ), .IFB94B817F0BC84EC0734110F6EDE475A (IB5B3486ECA0F911FF5D92A37ECF53B4A ), .I512A575E055CF9235066DBE4051242CB
(I0B5E80731173820DE30A1D6C548B918B ), .I391BF6A9C9F2ABEEA227F0E1F3F50A4F (I8A848F283F0A33BC04B5173E5E3FE015 ), .IF0D7F78B99E50997A728E3731A197225
(I0069A39965C0330678D64B612F60F78D ), .I9606837003EFA36A64A97C352D3D89A3 (I30A298A8327798F01C20DDAD6A556FB3 ), .I4C1994114E1C49B9376320858F4E71F9
(I4EB1044CFC38A54424DBAA59B9641ED6 ), .I2CB8399B2A61CDA9DB269D3567018E65 (IC920957C9C4BA12361B2EB75CD52EA74 ), .I46C5269B9FB24EF04CE2CC341C288EC7
(I46C5269B9FB24EF04CE2CC341C288EC7 ), .I3C9AD458B89B2FAABD743BF4E13BF421 (I3C9AD458B89B2FAABD743BF4E13BF421 ), .I73ABD5619A9FB885445AC1E288EAF7F8
(2), .IBDE0431C8F903800F409661F4F56FD80 (IB26EBF559CA483EACBAD1BCA4C580AF2 ) ) ID078DD71CF03D7FD68F95041DED5D5CE
( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ),
.ICB680FEAB46B6D635CD9DD6BB49A6A20 (IAA6C398FE19CA194DA9436764C94079A ), .I8FF768DAF4C56D1B2D217B2C02B6D4EC (I6375C05D4E0F58631C8731FD2B26A7F6 ),
.I9E5E6E86745F53F982BC3862031A206B (ID25293C6DC5461B1A3E61F7A7614A6D8 ), .I3AD72E1D6C16169DB8A27F1681293009 (I7E0B227F296E6A7FA770C68AB70324DD ),
.I0DE44F162EF92573C5DE1249527F6E9D (I1187CE134A1A3347BF94366BE4D44B3F ), .I2E9CC9AFC2E4742F852CB037CFC7E0A1 (I0C7C3FDEC159F63C155144A19841E5BC ),
.I8B1798242C3B0E655181D0D365813614 (I8B1798242C3B0E655181D0D365813614 ), .IE145222FDBDC80109E12FA72D3D3C655 (IE145222FDBDC80109E12FA72D3D3C655 ),
.ID43AC1009727D128F1C5DFE4640CA5AB (ID43AC1009727D128F1C5DFE4640CA5AB ), .IB610431939CB8180EAC2403672BAF58D (IB610431939CB8180EAC2403672BAF58D ),
.I3C7A9FA839F554D8898020C4831479E2 (IC7DB18773990D347CEF55E672D6B2C05 ), .I74A0936EE8FD1443A2C6745A4F3F6B5E (I39A06B46F4E1C11EE4BFB781E3B4F32A ),
.I369BA2FFB5D41DF25F9BC3AB126D6607 (I369BA2FFB5D41DF25F9BC3AB126D6607 ), .I1C0271AD5E8E9E9164909E468AD0B212 (IB4CA57E47B085EE5925036D5223A4598 ),
.I6EC1BE4B18EC6AA3D88A5D45B614565E (I6EC1BE4B18EC6AA3D88A5D45B614565E [2]), .I56148DDDF284443347FFCF4F9C3BE61A (I81BF37FCB51B492DCA857F28ABD8D76E [2]),
.I24C403550AE065D7D1B7266142886226 (I24C403550AE065D7D1B7266142886226 ), .I438B8BD876741F9B46EB770E92F808B7 (I438B8BD876741F9B46EB770E92F808B7 [11:0]),
.I5FE75BE614D4F52DB327549B36203350 (I74CF4D6FE5B30BB30E40AFCA2A08A220 [2]), .I3D6C771D05CA1A769E61302C086494B8 (I3D6C771D05CA1A769E61302C086494B8 ),
.I357B3043EDACE3EBECE8F54D79B9F90A (I357B3043EDACE3EBECE8F54D79B9F90A ), .I0AAD559CF33A5CBA597990658774FEB3 (I0AAD559CF33A5CBA597990658774FEB3 ),
.I923204A95D8CBB206587CF32BEDCF4EF (I923204A95D8CBB206587CF32BEDCF4EF ), .ICF9D8FD31DFC7D20DAF939C6D75F1518 (ICF9D8FD31DFC7D20DAF939C6D75F1518 [2]),
.IDF550B17734BF16B7E410B19BB31E276 (IB1AAAED8469CADFA3AB4BF806A8466B6 ), .I8ED9B9C1D9F58C5D06A9443AD901E8C6 (IA6774F4F4F3AF83C6A9E233DB00F89A0 ),
.IA976D63BEECA80DCE31365CF56EC0248 (IFFF50035216FD68A74F8164F0EE74689 ), .I5E3CE5AF5C34D232BFB139B63D9912B4 (IF9A16909C25386742335A246DEDE12E8 ),
.IBEF3E5F9395E2C7822AE03D6461DEBBB (I5078F81AE0F5DCD4CC2ABEE2CEF9C827 ), .I7E6CFD6A7DCAB9CD2188D044C7D716A6 (IB55475954FE95F83F22B1C2FB76FAEC7 ),
.I3A34691662384260F0524DD7F650E75A (I31980ABC07D19BA89784085C7754DE42 ), .IC2F58AB5028C1D2C53C6EF47A4975D0A (IE1F9397E899B4E938A0D54FC51445C13 ),
.I112E0A79129A8BC6DD4C13647C31F8A0 (IDE0F2D42601304C0E0CCD60778B3938F ), .IE4B6DD43E04940631EF58BA04EA58997 (IACF97B89AE62537A26788BDFCE846ED1 [2]),
.I3A095084CDFDFA56A0E67616A78D3B25 (I01D4C6B20466D26621C6DA5816817455 [2]), .I81CD7F184DF8D58A1F2324E975A6816C (I46A701488EBE724B47736C3C7A47A876 [2]),
.I83C4A4200EB2B3F6766D338284ECAAAF (IFE63F76C2A46B87271596BE8D0FFD21A [2]), .I42A419EB6EB8D11234AC3B2BCA0AE593 (IAF2A92B584FD036A9F751EB8F3FA7ACD ),
.IA41AC3CC6BC050DDC172724AB311315B (I5CF35907FA895D81AAC1AAFED86DBE1F ), .I31CF69FF368B36B4D6612DF16B3ABC6B (I21EE6CA5EBC86B66AC5EE8AF763FB838 [2]),
.IFE4A8CBA73734C6F0F0A078027E053D4 (IFFB9EED620356BDFB94697DB3606174F ), .ID7A2A8B1E9D92B60194D5FAFAAB15208 (I2C072E656BFCADF4877B42244D6D2307 ),
.IF274FAF97F5BACD693913BB418717A9D (IB96A9322FAF5941DF70737CA69F152A3 ), .ID95C13E7EE1CFE6A8743FF9E62C25873 (I5B92AFCE2F6F881BA10FA726B18BB692 ),
.IC58E411F24D810EF60A7B8638ABCC0BB (I60F6B756CD1062B40CC02E1438F28711 ), .I89CFFA73C7546481B72B0FB06D799AEE (I746F8C8440813F740701D80A6F08674F ),
.I270ED686C2EF2C1C8B5B55EC4A5AAE84 (I9625E96E33563830A2A0ED7263124B10 ), .ID5CCD4858CB5CC1B2EDEC682C7DE5AAD (I1B43D1CE930FCA067FA31726F2C15FEE ),
.I7D901091F9E0741061C75B54467D48A0 (I697639B04C0F4B6F9764F8122329FB7C ) ); else begin assign ICF9D8FD31DFC7D20DAF939C6D75F1518 [2]
= 1'b0; assign IACF97B89AE62537A26788BDFCE846ED1 [2] = 1'b0; assign I01D4C6B20466D26621C6DA5816817455 [2] = 1'b0;
assign I46A701488EBE724B47736C3C7A47A876 [2] = 1'b0; assign IFE63F76C2A46B87271596BE8D0FFD21A [2] = 1'b0; assign
I21EE6CA5EBC86B66AC5EE8AF763FB838 [2] = 1'b0; assign IB1AAAED8469CADFA3AB4BF806A8466B6 = 1'b0; assign IA6774F4F4F3AF83C6A9E233DB00F89A0
= 1'b0; assign IFFF50035216FD68A74F8164F0EE74689 = 1'b0; assign IF9A16909C25386742335A246DEDE12E8 = 1'b0; assign
I5078F81AE0F5DCD4CC2ABEE2CEF9C827 = 1'b0; assign IB55475954FE95F83F22B1C2FB76FAEC7 = 1'b0; assign I31980ABC07D19BA89784085C7754DE42
= 1'b0; assign IE1F9397E899B4E938A0D54FC51445C13 = 1'b0; assign IDE0F2D42601304C0E0CCD60778B3938F = 3'b0; assign
IAF2A92B584FD036A9F751EB8F3FA7ACD = 3'b0; assign I5CF35907FA895D81AAC1AAFED86DBE1F = 3'b0; assign IFFB9EED620356BDFB94697DB3606174F
= 32'b0; assign I2C072E656BFCADF4877B42244D6D2307 = 1'b0; assign IB96A9322FAF5941DF70737CA69F152A3 = 1'b0; assign
I5B92AFCE2F6F881BA10FA726B18BB692 = 1'b0; assign I60F6B756CD1062B40CC02E1438F28711 = 11'b0; assign I746F8C8440813F740701D80A6F08674F
= 1'b0; assign I9625E96E33563830A2A0ED7263124B10 = 1'b0; assign I1B43D1CE930FCA067FA31726F2C15FEE = 1'b0; assign
I697639B04C0F4B6F9764F8122329FB7C = 32'b0; end endgenerate  generate if (IFA272F301A5935EE15CB134524665363 ) I2296FC491415818D18357D6C2D700C14
# ( .IFC1FF746397E6A576E9FEB281890A248 (IB231E22D146559D11318B25AE0BA8C7A ), .IAF1DF965ED0D670C125D16FDF91B875B
(I7377F8B5325C7EE7D12D8B4B6A18183F ), .IB7B379BA36F36F0638F4F33C7598CC85 (I17C1305CE886D24D942A2A62C4DB3617 ), .ID9DCCEB6B5B42C479CB9D2B3C992035D
(ID926607BDA4008824BC8A9A1B67C04B7 ), .I251C6E5612F7B344EC3156CB9A93BE5B (IE4511A2FC6AD3FBAEAADD1EF75F0B773 ), .ID7A688D3DA9A2C539FE87FC8998248CB
(I0B29563399BE9E04B2FE3DE714C7DCE6 ), .I96DBC3D130FB2B57DFB76E3E87DF89D2 (I698853A251199BE8A5753717E876DA52 ), .I87B53E44EDBDCDA1796FB105323D3B17
(IA3BC4D015F529FD7E88E1370A882D0DF ), .IF9554E0938E353BDC05ABE0C628E3BE9 (I3463AC2A02018CF2288043A9C3E47A4F ), .I37C708634F442A3B0568DA0BB576511F
(IFDC235A84B81F7EB6EA5B1ED1F71197F ), .I7B125DA60401B7C86EB027E9E9262847 (IF0C0D849F42A4C05A7BF373811D5F5F5 ), .I8BEE88809FA5712893BC59FF0E17ADB2
(I59B19D300B55C10DB1B10364E9E59201 ), .I7DF5A90920A562D09AA22D2DFA657124 (IB1CD9FD007D322042A1087AC76B782B4 ), .I0243B4A4E84E0712929C806F438E6AA9
(I6A959CC2CFE148A0D8579A1CEE0C6699 ), .I7050B96C0C45A812BBFC45C2A30F272C (I1953E43D30396B1EDBD48DAD13C6A240 ), .IB7C70D5D7B0DDF146F4D402BEE6F6FA6
(IC02B62ACA36F1FEBB031FE435BA48A9A ), .I1CBD8B214B4765FBC7FA828F0C62BC94 (IAE6C36DBDB6FF8E962D96D8F1FB95CC1 ), .I677BE3663880CBE6E5AE2C431F3FDD4D
(I82E91D4ACF151209B3234E6F867049F1 ), .I1CF1EE9FA60C0CDB15DD404CC8A269E5 (I9806BFEA675277E4572CB4FD0C9C0D8C ), .I34F020684BFF4B1EAA406E693751B71D
(I802B81175874E1E34C3E4EE6C7F0B969 ), .IFB94B817F0BC84EC0734110F6EDE475A (I00773A8B25BA28541FF04BC530185E7F ), .I512A575E055CF9235066DBE4051242CB
(IB2267C4E34709B9CE9D697340B9DA12F ), .I391BF6A9C9F2ABEEA227F0E1F3F50A4F (I37AC0331E13434E399C90A5408FB09E2 ), .IF0D7F78B99E50997A728E3731A197225
(IC69BEB80DB094A65F3DFB0265F8616DE ), .I9606837003EFA36A64A97C352D3D89A3 (I6C4A37BD8E4A0A1D9639A3FA64D5F8C3 ), .I4C1994114E1C49B9376320858F4E71F9
(ID969B30E2BD8213873A2D19FFDEF204A ), .I2CB8399B2A61CDA9DB269D3567018E65 (IC3F1AF003F5E2257563771F88647B5FF ), .I46C5269B9FB24EF04CE2CC341C288EC7
(I46C5269B9FB24EF04CE2CC341C288EC7 ), .I3C9AD458B89B2FAABD743BF4E13BF421 (I3C9AD458B89B2FAABD743BF4E13BF421 ), .I73ABD5619A9FB885445AC1E288EAF7F8
(3), .IBDE0431C8F903800F409661F4F56FD80 (IB26EBF559CA483EACBAD1BCA4C580AF2 ) ) ICD3794690C7B631F413EC5D0D0043A96
( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ),
.ICB680FEAB46B6D635CD9DD6BB49A6A20 (IF0C365E1D4BC8B2941DE257EF66C8FE4 ), .I8FF768DAF4C56D1B2D217B2C02B6D4EC (I1646E818A90159BC4FF7AA119272C460 ),
.I9E5E6E86745F53F982BC3862031A206B (I05AD49E3884F0E62FA36DCFB88E5C22E ), .I3AD72E1D6C16169DB8A27F1681293009 (I348CE8EA5A014339F820FDCAFC214867 ),
.I0DE44F162EF92573C5DE1249527F6E9D (ICF2AC2986B60A3FD41ECFB74C4756D10 ), .I2E9CC9AFC2E4742F852CB037CFC7E0A1 (I13B899B342E8552CACED9E20E0F5FD83 ),
.I8B1798242C3B0E655181D0D365813614 (I8B1798242C3B0E655181D0D365813614 ), .IE145222FDBDC80109E12FA72D3D3C655 (IE145222FDBDC80109E12FA72D3D3C655 ),
.ID43AC1009727D128F1C5DFE4640CA5AB (ID43AC1009727D128F1C5DFE4640CA5AB ), .IB610431939CB8180EAC2403672BAF58D (IB610431939CB8180EAC2403672BAF58D ),
.I3C7A9FA839F554D8898020C4831479E2 (IC7DB18773990D347CEF55E672D6B2C05 ), .I74A0936EE8FD1443A2C6745A4F3F6B5E (I39A06B46F4E1C11EE4BFB781E3B4F32A ),
.I369BA2FFB5D41DF25F9BC3AB126D6607 (I369BA2FFB5D41DF25F9BC3AB126D6607 ), .I1C0271AD5E8E9E9164909E468AD0B212 (I2F92739468FA7128C93936C8511AA228 ),
.I6EC1BE4B18EC6AA3D88A5D45B614565E (I6EC1BE4B18EC6AA3D88A5D45B614565E [3]), .I56148DDDF284443347FFCF4F9C3BE61A (I81BF37FCB51B492DCA857F28ABD8D76E [3]),
.I24C403550AE065D7D1B7266142886226 (I24C403550AE065D7D1B7266142886226 ), .I438B8BD876741F9B46EB770E92F808B7 (I438B8BD876741F9B46EB770E92F808B7 [11:0]),
.I5FE75BE614D4F52DB327549B36203350 (I74CF4D6FE5B30BB30E40AFCA2A08A220 [3]), .I3D6C771D05CA1A769E61302C086494B8 (I3D6C771D05CA1A769E61302C086494B8 ),
.I357B3043EDACE3EBECE8F54D79B9F90A (I357B3043EDACE3EBECE8F54D79B9F90A ), .I0AAD559CF33A5CBA597990658774FEB3 (I0AAD559CF33A5CBA597990658774FEB3 ),
.I923204A95D8CBB206587CF32BEDCF4EF (I923204A95D8CBB206587CF32BEDCF4EF ), .ICF9D8FD31DFC7D20DAF939C6D75F1518 (ICF9D8FD31DFC7D20DAF939C6D75F1518 [3]),
.IDF550B17734BF16B7E410B19BB31E276 (I1E1A1AD224EE52C02213B0661856A826 ), .I8ED9B9C1D9F58C5D06A9443AD901E8C6 (IDBF2DE7607B69A821EF14BD65A75A2DC ),
.IA976D63BEECA80DCE31365CF56EC0248 (IB35E0CDEF8AAA93EF9B0047DE75BCDB1 ), .I5E3CE5AF5C34D232BFB139B63D9912B4 (IC5663A92559813188629C72D2AF75E2B ),
.IBEF3E5F9395E2C7822AE03D6461DEBBB (IB7ADE2C78FA2211545637C290CFB45CB ), .I7E6CFD6A7DCAB9CD2188D044C7D716A6 (I38BDB4EBCC779338E7AF863601C4853E ),
.I3A34691662384260F0524DD7F650E75A (ICD34F2C7357A369358E7CFBC3D425106 ), .IC2F58AB5028C1D2C53C6EF47A4975D0A (I081CFEF0428EFE96BD06A8F2EE9DC2CD ),
.I112E0A79129A8BC6DD4C13647C31F8A0 (ID34187ADCB71E296DE727A7573E76A15 ), .IE4B6DD43E04940631EF58BA04EA58997 (IACF97B89AE62537A26788BDFCE846ED1 [3]),
.I3A095084CDFDFA56A0E67616A78D3B25 (I01D4C6B20466D26621C6DA5816817455 [3]), .I81CD7F184DF8D58A1F2324E975A6816C (I46A701488EBE724B47736C3C7A47A876 [3]),
.I83C4A4200EB2B3F6766D338284ECAAAF (IFE63F76C2A46B87271596BE8D0FFD21A [3]), .I42A419EB6EB8D11234AC3B2BCA0AE593 (I5B6B84BEB62496031A951D18F8043152 ),
.IA41AC3CC6BC050DDC172724AB311315B (IC21D6CA5169E489082288A960FB9DDFE ), .I31CF69FF368B36B4D6612DF16B3ABC6B (I21EE6CA5EBC86B66AC5EE8AF763FB838 [3]),
.IFE4A8CBA73734C6F0F0A078027E053D4 (I0D8A716B0016AFE64E7F7977A80A253A ), .ID7A2A8B1E9D92B60194D5FAFAAB15208 (IAEFBAA4728FB6854C056C8E4C0691B3D ),
.IF274FAF97F5BACD693913BB418717A9D (I1DC328E1B03775141AFCFBB60C78CDC0 ), .ID95C13E7EE1CFE6A8743FF9E62C25873 (I3ABE7E8A0A3ADCF18D9C06A84D938210 ),
.IC58E411F24D810EF60A7B8638ABCC0BB (I6DA6F40C5003D56BA074AD254DFE4B48 ), .I89CFFA73C7546481B72B0FB06D799AEE (I55D773F0648256E2B67F14A58A7AE480 ),
.I270ED686C2EF2C1C8B5B55EC4A5AAE84 (I0F56078C1F80B8234A46BCE05F251A14 ), .ID5CCD4858CB5CC1B2EDEC682C7DE5AAD (IA37321C9DB7C6279A1BBB82432DD22B2 ),
.I7D901091F9E0741061C75B54467D48A0 (I3C0E217327A8665923FDC969639C89C7 ) ); else begin assign ICF9D8FD31DFC7D20DAF939C6D75F1518 [3]
= 1'b0; assign IACF97B89AE62537A26788BDFCE846ED1 [3] = 1'b0; assign I01D4C6B20466D26621C6DA5816817455 [3] = 1'b0;
assign I46A701488EBE724B47736C3C7A47A876 [3] = 1'b0; assign IFE63F76C2A46B87271596BE8D0FFD21A [3] = 1'b0; assign
I21EE6CA5EBC86B66AC5EE8AF763FB838 [3] = 1'b0; assign I1E1A1AD224EE52C02213B0661856A826 = 1'b0; assign IDBF2DE7607B69A821EF14BD65A75A2DC
= 1'b0; assign IB35E0CDEF8AAA93EF9B0047DE75BCDB1 = 1'b0; assign IC5663A92559813188629C72D2AF75E2B = 1'b0; assign
IB7ADE2C78FA2211545637C290CFB45CB = 1'b0; assign I38BDB4EBCC779338E7AF863601C4853E = 1'b0; assign ICD34F2C7357A369358E7CFBC3D425106
= 1'b0; assign I081CFEF0428EFE96BD06A8F2EE9DC2CD = 1'b0; assign ID34187ADCB71E296DE727A7573E76A15 = 3'b0; assign
I5B6B84BEB62496031A951D18F8043152 = 3'b0; assign IC21D6CA5169E489082288A960FB9DDFE = 3'b0; assign I0D8A716B0016AFE64E7F7977A80A253A
= 32'b0; assign IAEFBAA4728FB6854C056C8E4C0691B3D = 1'b0; assign I1DC328E1B03775141AFCFBB60C78CDC0 = 1'b0; assign
I3ABE7E8A0A3ADCF18D9C06A84D938210 = 1'b0; assign I6DA6F40C5003D56BA074AD254DFE4B48 = 11'b0; assign I55D773F0648256E2B67F14A58A7AE480
= 1'b0; assign I0F56078C1F80B8234A46BCE05F251A14 = 1'b0; assign IA37321C9DB7C6279A1BBB82432DD22B2 = 1'b0; assign
I3C0E217327A8665923FDC969639C89C7 = 32'b0; end endgenerate  generate if (IE690B7723F136DA02896C0728DDADB49 ) I2296FC491415818D18357D6C2D700C14
# ( .IFC1FF746397E6A576E9FEB281890A248 (I21752C34E9BF9458DB0D20BA11A8898B ), .IAF1DF965ED0D670C125D16FDF91B875B
(IBFD9199C154D56895B673A496CF82DA3 ), .IB7B379BA36F36F0638F4F33C7598CC85 (I900E9757930519C7865CA2247E6CC23A ), .ID9DCCEB6B5B42C479CB9D2B3C992035D
(IFA7D0D435AE6BBF59445626F82B8B26E ), .I251C6E5612F7B344EC3156CB9A93BE5B (IA794CD2FEB24AB956EC1914852D2E7D5 ), .ID7A688D3DA9A2C539FE87FC8998248CB
(IAED1399D2D60713A0101069DD427D0A0 ), .I96DBC3D130FB2B57DFB76E3E87DF89D2 (I72E6ED810779933C7E2125FC345DEC0B ), .I87B53E44EDBDCDA1796FB105323D3B17
(I3C7842C10567F9851F14519598E7EE93 ), .IF9554E0938E353BDC05ABE0C628E3BE9 (I1DE5880AD46DABF7282A3FF245F71602 ), .I37C708634F442A3B0568DA0BB576511F
(I7747208BC7A624CD71D5BB421E9EE4A4 ), .I7B125DA60401B7C86EB027E9E9262847 (I4103D81EBFB4946FA8F9593A8B7DE5C8 ), .I8BEE88809FA5712893BC59FF0E17ADB2
(I858B464778E6994385995C3205FB37B0 ), .I7DF5A90920A562D09AA22D2DFA657124 (I785E686713BEF380843045D4DB00E51C ), .I0243B4A4E84E0712929C806F438E6AA9
(IABD30C53E56587015015FE5F556929D7 ), .I7050B96C0C45A812BBFC45C2A30F272C (IABB4198D13BE4058E856EBC11D8D6565 ), .IB7C70D5D7B0DDF146F4D402BEE6F6FA6
(I0405497FA63FB5AA449F0C813D8E8F89 ), .I1CBD8B214B4765FBC7FA828F0C62BC94 (I6F86DD61D81AE7AE015C945BA5CF8828 ), .I677BE3663880CBE6E5AE2C431F3FDD4D
(I69C4352219E15BD98C0B6A7428BAB037 ), .I1CF1EE9FA60C0CDB15DD404CC8A269E5 (I68ED8551754B5BAA65EB2F191A697C4B ), .I34F020684BFF4B1EAA406E693751B71D
(ICE0C22941CF3ECFDB4B47576E4E4A06E ), .IFB94B817F0BC84EC0734110F6EDE475A (I262F500CDAF1182E64A895FA5F58D006 ), .I512A575E055CF9235066DBE4051242CB
(ID88F3DF54AD4CA3D33C94EC1E1B5BB01 ), .I391BF6A9C9F2ABEEA227F0E1F3F50A4F (I8F019158F18BA70FE5953E859D4BA891 ), .IF0D7F78B99E50997A728E3731A197225
(I4046611EA3EEF60ACE26738C818FDBA2 ), .I9606837003EFA36A64A97C352D3D89A3 (I78E815C8C6F11755E08393F339C5E874 ), .I4C1994114E1C49B9376320858F4E71F9
(IC377F0EF36016932385B3B0988B91B0F ), .I2CB8399B2A61CDA9DB269D3567018E65 (IBDEA2513680CC11B2E5E42FB17332F70 ), .I46C5269B9FB24EF04CE2CC341C288EC7
(I46C5269B9FB24EF04CE2CC341C288EC7 ), .I3C9AD458B89B2FAABD743BF4E13BF421 (I3C9AD458B89B2FAABD743BF4E13BF421 ), .I73ABD5619A9FB885445AC1E288EAF7F8
(4), .IBDE0431C8F903800F409661F4F56FD80 (IB26EBF559CA483EACBAD1BCA4C580AF2 ) ) I163D5B15D15A52B858B1A6A5B84A887B
( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ),
.ICB680FEAB46B6D635CD9DD6BB49A6A20 (I068B3206EC02BBE1225E3FD649DCAC3E ), .I8FF768DAF4C56D1B2D217B2C02B6D4EC (I15D8A1D8934ABE732F753BC8A130129E ),
.I9E5E6E86745F53F982BC3862031A206B (IFE8F569C18FBA7444D4832F2CB5D2D69 ), .I3AD72E1D6C16169DB8A27F1681293009 (I51FF9F99E3F92A151FD3D6BBAAC89FB6 ),
.I0DE44F162EF92573C5DE1249527F6E9D (IA4118298EF0A9C92D5D3ECB07C8AE533 ), .I2E9CC9AFC2E4742F852CB037CFC7E0A1 (I7D032A1E448C6F22898894E594BF2DD3 ),
.I8B1798242C3B0E655181D0D365813614 (I8B1798242C3B0E655181D0D365813614 ), .IE145222FDBDC80109E12FA72D3D3C655 (IE145222FDBDC80109E12FA72D3D3C655 ),
.ID43AC1009727D128F1C5DFE4640CA5AB (ID43AC1009727D128F1C5DFE4640CA5AB ), .IB610431939CB8180EAC2403672BAF58D (IB610431939CB8180EAC2403672BAF58D ),
.I3C7A9FA839F554D8898020C4831479E2 (IC7DB18773990D347CEF55E672D6B2C05 ), .I74A0936EE8FD1443A2C6745A4F3F6B5E (I39A06B46F4E1C11EE4BFB781E3B4F32A ),
.I369BA2FFB5D41DF25F9BC3AB126D6607 (I369BA2FFB5D41DF25F9BC3AB126D6607 ), .I1C0271AD5E8E9E9164909E468AD0B212 (I25DCCEF37BE2FCC042C00B81ABCA449F ),
.I6EC1BE4B18EC6AA3D88A5D45B614565E (I6EC1BE4B18EC6AA3D88A5D45B614565E [4]), .I56148DDDF284443347FFCF4F9C3BE61A (I81BF37FCB51B492DCA857F28ABD8D76E [4]),
.I24C403550AE065D7D1B7266142886226 (I24C403550AE065D7D1B7266142886226 ), .I438B8BD876741F9B46EB770E92F808B7 (I438B8BD876741F9B46EB770E92F808B7 [11:0]),
.I5FE75BE614D4F52DB327549B36203350 (I74CF4D6FE5B30BB30E40AFCA2A08A220 [4]), .I3D6C771D05CA1A769E61302C086494B8 (I3D6C771D05CA1A769E61302C086494B8 ),
.I357B3043EDACE3EBECE8F54D79B9F90A (I357B3043EDACE3EBECE8F54D79B9F90A ), .I0AAD559CF33A5CBA597990658774FEB3 (I0AAD559CF33A5CBA597990658774FEB3 ),
.I923204A95D8CBB206587CF32BEDCF4EF (I923204A95D8CBB206587CF32BEDCF4EF ), .ICF9D8FD31DFC7D20DAF939C6D75F1518 (ICF9D8FD31DFC7D20DAF939C6D75F1518 [4]),
.IDF550B17734BF16B7E410B19BB31E276 (I22F7EBEFD72C22C64DB546CE211C3C33 ), .I8ED9B9C1D9F58C5D06A9443AD901E8C6 (I7DA4C0DA5661A2191D932C4F426DE5F4 ),
.IA976D63BEECA80DCE31365CF56EC0248 (I17B065631E7403BD94AABA998687E920 ), .I5E3CE5AF5C34D232BFB139B63D9912B4 (I2D58D8090233025B63B11977CCF7A6FB ),
.IBEF3E5F9395E2C7822AE03D6461DEBBB (I79527CA6375BFC9B46B48DEFE32DEEAA ), .I7E6CFD6A7DCAB9CD2188D044C7D716A6 (I270710745C28824E285C2E05FB618D27 ),
.I3A34691662384260F0524DD7F650E75A (I765A5C6CB6D2AE7496EF2BE962529E09 ), .IC2F58AB5028C1D2C53C6EF47A4975D0A (I9C559D18449178998B7475813A7D0CBB ),
.I112E0A79129A8BC6DD4C13647C31F8A0 (I7B62DE436B5B4C0A20CC4FE1E5D6F91D ), .IE4B6DD43E04940631EF58BA04EA58997 (IACF97B89AE62537A26788BDFCE846ED1 [4]),
.I3A095084CDFDFA56A0E67616A78D3B25 (I01D4C6B20466D26621C6DA5816817455 [4]), .I81CD7F184DF8D58A1F2324E975A6816C (I46A701488EBE724B47736C3C7A47A876 [4]),
.I83C4A4200EB2B3F6766D338284ECAAAF (IFE63F76C2A46B87271596BE8D0FFD21A [4]), .I42A419EB6EB8D11234AC3B2BCA0AE593 (I56408FACA355983EAB06294FBFDA5C73 ),
.IA41AC3CC6BC050DDC172724AB311315B (IDAF814B27DE872458FE905492366EC1F ), .I31CF69FF368B36B4D6612DF16B3ABC6B (I21EE6CA5EBC86B66AC5EE8AF763FB838 [4]),
.IFE4A8CBA73734C6F0F0A078027E053D4 (I88DEF602C28E2AE7FCFC75761E9DF8F6 ), .ID7A2A8B1E9D92B60194D5FAFAAB15208 (I6434FE6B1DB9B4DCDB82F1E568D8A5AD ),
.IF274FAF97F5BACD693913BB418717A9D (IF76FEAB2FA7E91BC33928D6B232B6040 ), .ID95C13E7EE1CFE6A8743FF9E62C25873 (IA3A543EBA3F35D293D9F9A372241FFB7 ),
.IC58E411F24D810EF60A7B8638ABCC0BB (I6913053E317EA8A5066057EFF8119A7D ), .I89CFFA73C7546481B72B0FB06D799AEE (I96F424D83A110B76A1E3957956BB0EEA ),
.I270ED686C2EF2C1C8B5B55EC4A5AAE84 (ID24D46A573CB38B617C5B4569142A8C0 ), .ID5CCD4858CB5CC1B2EDEC682C7DE5AAD (I097D8CB350937ECACE8C02CAB12CF7F5 ),
.I7D901091F9E0741061C75B54467D48A0 (ID04E1BCD61D6D921C4E551FD2CE92041 ) ); else begin assign ICF9D8FD31DFC7D20DAF939C6D75F1518 [4]
= 1'b0; assign IACF97B89AE62537A26788BDFCE846ED1 [4] = 1'b0; assign I01D4C6B20466D26621C6DA5816817455 [4] = 1'b0;
assign I46A701488EBE724B47736C3C7A47A876 [4] = 1'b0; assign IFE63F76C2A46B87271596BE8D0FFD21A [4] = 1'b0; assign
I21EE6CA5EBC86B66AC5EE8AF763FB838 [4] = 1'b0; assign I22F7EBEFD72C22C64DB546CE211C3C33 = 1'b0; assign I7DA4C0DA5661A2191D932C4F426DE5F4
= 1'b0; assign I17B065631E7403BD94AABA998687E920 = 1'b0; assign I2D58D8090233025B63B11977CCF7A6FB = 1'b0; assign
I79527CA6375BFC9B46B48DEFE32DEEAA = 1'b0; assign I270710745C28824E285C2E05FB618D27 = 1'b0; assign I765A5C6CB6D2AE7496EF2BE962529E09
= 1'b0; assign I9C559D18449178998B7475813A7D0CBB = 1'b0; assign I7B62DE436B5B4C0A20CC4FE1E5D6F91D = 3'b0; assign
I56408FACA355983EAB06294FBFDA5C73 = 3'b0; assign IDAF814B27DE872458FE905492366EC1F = 3'b0; assign I88DEF602C28E2AE7FCFC75761E9DF8F6
= 32'b0; assign I6434FE6B1DB9B4DCDB82F1E568D8A5AD = 1'b0; assign IF76FEAB2FA7E91BC33928D6B232B6040 = 1'b0; assign
IA3A543EBA3F35D293D9F9A372241FFB7 = 1'b0; assign I6913053E317EA8A5066057EFF8119A7D = 11'b0; assign I96F424D83A110B76A1E3957956BB0EEA
= 1'b0; assign ID24D46A573CB38B617C5B4569142A8C0 = 1'b0; assign I097D8CB350937ECACE8C02CAB12CF7F5 = 1'b0; assign
ID04E1BCD61D6D921C4E551FD2CE92041 = 32'b0; end endgenerate  generate if (I55BE27080C370AF723A4FE096014E875 ) I2296FC491415818D18357D6C2D700C14
# ( .IFC1FF746397E6A576E9FEB281890A248 (IDC77C35F0E8480627E0F64F68D8A39ED ), .IAF1DF965ED0D670C125D16FDF91B875B
(I110F59F054A1064BFB27909E2370F028 ), .IB7B379BA36F36F0638F4F33C7598CC85 (IED76B05540143124D123636B36A006DA ), .ID9DCCEB6B5B42C479CB9D2B3C992035D
(I96B06C30CEFF410BD39B69C003D2AC2B ), .I251C6E5612F7B344EC3156CB9A93BE5B (I2050954950618B2F390C43E2A3A4A814 ), .ID7A688D3DA9A2C539FE87FC8998248CB
(I3F39386711BA6D94D8C7A1C5710875D6 ), .I96DBC3D130FB2B57DFB76E3E87DF89D2 (I3011FF9154FC5D6F394688805C3D9B33 ), .I87B53E44EDBDCDA1796FB105323D3B17
(I08E7BC06415AD0F55BE9EFFEB79B0315 ), .IF9554E0938E353BDC05ABE0C628E3BE9 (IB069DEA93E56D26CAB0E5B9C9E284CDE ), .I37C708634F442A3B0568DA0BB576511F
(I5F80A9459505144CBBE328F0713782CC ), .I7B125DA60401B7C86EB027E9E9262847 (IC88E0007329C31C00B55FD745AAD6590 ), .I8BEE88809FA5712893BC59FF0E17ADB2
(I102247373FC0AC7EA52B3EFB2A5CC280 ), .I7DF5A90920A562D09AA22D2DFA657124 (I750129419895285C7D4ABEB3C2FEEE71 ), .I0243B4A4E84E0712929C806F438E6AA9
(I2CFDEF4EE4DDBFD88BE646118F3E6FE2 ), .I7050B96C0C45A812BBFC45C2A30F272C (ID42754EA33A6C985294D5AD602396DA3 ), .IB7C70D5D7B0DDF146F4D402BEE6F6FA6
(I6FBC4AA1ED36E030778F1A24E9C9B2E4 ), .I1CBD8B214B4765FBC7FA828F0C62BC94 (I15A258E402E001F63FAB5BE8DF569399 ), .I677BE3663880CBE6E5AE2C431F3FDD4D
(IA2FE22B25B2F0C96B10399B2FB4B7C81 ), .I1CF1EE9FA60C0CDB15DD404CC8A269E5 (I36E46FAD7B2BA4DF9270A70F4921CC43 ), .I34F020684BFF4B1EAA406E693751B71D
(I0500A389ECC6C6D86EA16632126031AD ), .IFB94B817F0BC84EC0734110F6EDE475A (IFF2CDD869828E984763A775FF1821810 ), .I512A575E055CF9235066DBE4051242CB
(I4A7FAB30233B5A9954B6B6AD08DCADAA ), .I391BF6A9C9F2ABEEA227F0E1F3F50A4F (IC7B583F6D8F8A6C3C62D45FA87D50A19 ), .IF0D7F78B99E50997A728E3731A197225
(IAE03DAE231BA40E8DD1C02D38068EF8A ), .I9606837003EFA36A64A97C352D3D89A3 (IB842E33563B3EE1795267FE015C7B1A0 ), .I4C1994114E1C49B9376320858F4E71F9
(I229F764F8E53B82969E0B6B9234098CF ), .I2CB8399B2A61CDA9DB269D3567018E65 (IA9807BAB69B1AFAF9739BF86D99A92C3 ), .I46C5269B9FB24EF04CE2CC341C288EC7
(I46C5269B9FB24EF04CE2CC341C288EC7 ), .I3C9AD458B89B2FAABD743BF4E13BF421 (I3C9AD458B89B2FAABD743BF4E13BF421 ), .I73ABD5619A9FB885445AC1E288EAF7F8
(5), .IBDE0431C8F903800F409661F4F56FD80 (IB26EBF559CA483EACBAD1BCA4C580AF2 ) ) I1C325276098F305EDD5A96B670ED7E4B
( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ),
.ICB680FEAB46B6D635CD9DD6BB49A6A20 (I67444F97CA6B95448FAFAE30BC1EA4A3 ), .I8FF768DAF4C56D1B2D217B2C02B6D4EC (ID449FF330193AAA4C7942F23F18CEF54 ),
.I9E5E6E86745F53F982BC3862031A206B (I3CABF30E4ECE3E02DF7BB2FAE8895026 ), .I3AD72E1D6C16169DB8A27F1681293009 (I46EAD98AAF05965858087C6CCDFEAFFD ),
.I0DE44F162EF92573C5DE1249527F6E9D (I1967BD95F38270D97B0A4B182C5D8F0E ), .I2E9CC9AFC2E4742F852CB037CFC7E0A1 (ICDB8224D569BB5A5B320A26E2B451BAC ),
.I8B1798242C3B0E655181D0D365813614 (I8B1798242C3B0E655181D0D365813614 ), .IE145222FDBDC80109E12FA72D3D3C655 (IE145222FDBDC80109E12FA72D3D3C655 ),
.ID43AC1009727D128F1C5DFE4640CA5AB (ID43AC1009727D128F1C5DFE4640CA5AB ), .IB610431939CB8180EAC2403672BAF58D (IB610431939CB8180EAC2403672BAF58D ),
.I3C7A9FA839F554D8898020C4831479E2 (IC7DB18773990D347CEF55E672D6B2C05 ), .I74A0936EE8FD1443A2C6745A4F3F6B5E (I39A06B46F4E1C11EE4BFB781E3B4F32A ),
.I369BA2FFB5D41DF25F9BC3AB126D6607 (I369BA2FFB5D41DF25F9BC3AB126D6607 ), .I1C0271AD5E8E9E9164909E468AD0B212 (I19381BD04F07A020B45A7EFE952EBD90 ),
.I6EC1BE4B18EC6AA3D88A5D45B614565E (I6EC1BE4B18EC6AA3D88A5D45B614565E [5]), .I56148DDDF284443347FFCF4F9C3BE61A (I81BF37FCB51B492DCA857F28ABD8D76E [5]),
.I24C403550AE065D7D1B7266142886226 (I24C403550AE065D7D1B7266142886226 ), .I438B8BD876741F9B46EB770E92F808B7 (I438B8BD876741F9B46EB770E92F808B7 [11:0]),
.I5FE75BE614D4F52DB327549B36203350 (I74CF4D6FE5B30BB30E40AFCA2A08A220 [5]), .I3D6C771D05CA1A769E61302C086494B8 (I3D6C771D05CA1A769E61302C086494B8 ),
.I357B3043EDACE3EBECE8F54D79B9F90A (I357B3043EDACE3EBECE8F54D79B9F90A ), .I0AAD559CF33A5CBA597990658774FEB3 (I0AAD559CF33A5CBA597990658774FEB3 ),
.I923204A95D8CBB206587CF32BEDCF4EF (I923204A95D8CBB206587CF32BEDCF4EF ), .ICF9D8FD31DFC7D20DAF939C6D75F1518 (ICF9D8FD31DFC7D20DAF939C6D75F1518 [5]),
.IDF550B17734BF16B7E410B19BB31E276 (I0ED491A5B7F42029CCB818A7A566A126 ), .I8ED9B9C1D9F58C5D06A9443AD901E8C6 (I64422991E0FA499CEA26156FB729091E ),
.IA976D63BEECA80DCE31365CF56EC0248 (I1C44B39C210FB0191DFBF4FF9B4EB5AC ), .I5E3CE5AF5C34D232BFB139B63D9912B4 (IC3DC126AC872E9080FFE257241E00572 ),
.IBEF3E5F9395E2C7822AE03D6461DEBBB (IBCCBF2F5A49A76D461A7479DA2813EA7 ), .I7E6CFD6A7DCAB9CD2188D044C7D716A6 (IFFE90484B4E519D0DD55AFC0D9379B2A ),
.I3A34691662384260F0524DD7F650E75A (I6FDDB4608592CC601F82E29CF03F58E2 ), .IC2F58AB5028C1D2C53C6EF47A4975D0A (IE6E0B2D716FF39D4E07D15E9EAAB04FC ),
.I112E0A79129A8BC6DD4C13647C31F8A0 (IA2F68AF483F09457F392B22939441F47 ), .IE4B6DD43E04940631EF58BA04EA58997 (IACF97B89AE62537A26788BDFCE846ED1 [5]),
.I3A095084CDFDFA56A0E67616A78D3B25 (I01D4C6B20466D26621C6DA5816817455 [5]), .I81CD7F184DF8D58A1F2324E975A6816C (I46A701488EBE724B47736C3C7A47A876 [5]),
.I83C4A4200EB2B3F6766D338284ECAAAF (IFE63F76C2A46B87271596BE8D0FFD21A [5]), .I42A419EB6EB8D11234AC3B2BCA0AE593 (I8238B208D31228316827652162FA0720 ),
.IA41AC3CC6BC050DDC172724AB311315B (I28192CB07D936DD6F915E872C9D77566 ), .I31CF69FF368B36B4D6612DF16B3ABC6B (I21EE6CA5EBC86B66AC5EE8AF763FB838 [5]),
.IFE4A8CBA73734C6F0F0A078027E053D4 (I98308209671212A3C88A9644B503FA02 ), .ID7A2A8B1E9D92B60194D5FAFAAB15208 (IB4C822D6BFAE40F12254437B18142B8A ),
.IF274FAF97F5BACD693913BB418717A9D (I30157CAB406F288B630EF42C05ACC134 ), .ID95C13E7EE1CFE6A8743FF9E62C25873 (I82635882370B55739EA7454635CE3A41 ),
.IC58E411F24D810EF60A7B8638ABCC0BB (IE38989B54E8F0643FD2DC5F4F7B5BCC6 ), .I89CFFA73C7546481B72B0FB06D799AEE (I42E863B8B97EAE3620723BFD560E96F6 ),
.I270ED686C2EF2C1C8B5B55EC4A5AAE84 (I5ADEE764CD8A8EACE17ED8F55EC633AC ), .ID5CCD4858CB5CC1B2EDEC682C7DE5AAD (I977D818DD621CC225F1001F838F63684 ),
.I7D901091F9E0741061C75B54467D48A0 (I56C985EEB74E064645781DE4618A62B0 ) ); else begin assign ICF9D8FD31DFC7D20DAF939C6D75F1518 [5]
= 1'b0; assign IACF97B89AE62537A26788BDFCE846ED1 [5] = 1'b0; assign I01D4C6B20466D26621C6DA5816817455 [5] = 1'b0;
assign I46A701488EBE724B47736C3C7A47A876 [5] = 1'b0; assign IFE63F76C2A46B87271596BE8D0FFD21A [5] = 1'b0; assign
I21EE6CA5EBC86B66AC5EE8AF763FB838 [5] = 1'b0; assign I0ED491A5B7F42029CCB818A7A566A126 = 1'b0; assign I64422991E0FA499CEA26156FB729091E
= 1'b0; assign I1C44B39C210FB0191DFBF4FF9B4EB5AC = 1'b0; assign IC3DC126AC872E9080FFE257241E00572 = 1'b0; assign
IBCCBF2F5A49A76D461A7479DA2813EA7 = 1'b0; assign IFFE90484B4E519D0DD55AFC0D9379B2A = 1'b0; assign I6FDDB4608592CC601F82E29CF03F58E2
= 1'b0; assign IE6E0B2D716FF39D4E07D15E9EAAB04FC = 1'b0; assign IA2F68AF483F09457F392B22939441F47 = 3'b0; assign
I8238B208D31228316827652162FA0720 = 3'b0; assign I28192CB07D936DD6F915E872C9D77566 = 3'b0; assign I98308209671212A3C88A9644B503FA02
= 32'b0; assign IB4C822D6BFAE40F12254437B18142B8A = 1'b0; assign I30157CAB406F288B630EF42C05ACC134 = 1'b0; assign
I82635882370B55739EA7454635CE3A41 = 1'b0; assign IE38989B54E8F0643FD2DC5F4F7B5BCC6 = 11'b0; assign I42E863B8B97EAE3620723BFD560E96F6
= 1'b0; assign I5ADEE764CD8A8EACE17ED8F55EC633AC = 1'b0; assign I977D818DD621CC225F1001F838F63684 = 1'b0; assign
I56C985EEB74E064645781DE4618A62B0 = 32'b0; end endgenerate  generate if (IB2560D175E4507798B84D6E659FD6373 ) I2296FC491415818D18357D6C2D700C14
# ( .IFC1FF746397E6A576E9FEB281890A248 (IF02D8DF664D45B9699745A4C477F4220 ), .IAF1DF965ED0D670C125D16FDF91B875B
(I553DE26948BD8999C232161660D3E8AF ), .IB7B379BA36F36F0638F4F33C7598CC85 (IB99020DD53AEEF55E5DA5BF15890E9A5 ), .ID9DCCEB6B5B42C479CB9D2B3C992035D
(I0108C021E74AB8DE1357A170111B08CF ), .I251C6E5612F7B344EC3156CB9A93BE5B (IDED06CF1ED1692C601F91B904599696F ), .ID7A688D3DA9A2C539FE87FC8998248CB
(I7926E122D54A321BCD3309E19D9A0183 ), .I96DBC3D130FB2B57DFB76E3E87DF89D2 (I48C74401BD4D3F04619117E263213AFA ), .I87B53E44EDBDCDA1796FB105323D3B17
(I40F4EF6A18605258D6F6893B593AA318 ), .IF9554E0938E353BDC05ABE0C628E3BE9 (IAB56F2CB5ED41158B5A0ABE2FD915084 ), .I37C708634F442A3B0568DA0BB576511F
(I11F59D9A3377C9C28FB84219B4A4E4DC ), .I7B125DA60401B7C86EB027E9E9262847 (I3BE4D977225B6255BC284FA193DD9241 ), .I8BEE88809FA5712893BC59FF0E17ADB2
(I6A49481E89496C888774F840785C0BA4 ), .I7DF5A90920A562D09AA22D2DFA657124 (IE19B87A06C26E07981B4C116F5E878F7 ), .I0243B4A4E84E0712929C806F438E6AA9
(IF587F6E4A635FC1DA01C698D24B80510 ), .I7050B96C0C45A812BBFC45C2A30F272C (IBF68DF087726DF134221B625725579B8 ), .IB7C70D5D7B0DDF146F4D402BEE6F6FA6
(I9F10A6A60E1AEDF0BC22B2ED2686E4C2 ), .I1CBD8B214B4765FBC7FA828F0C62BC94 (I10394C1F82392903C22C104CEC600C4E ), .I677BE3663880CBE6E5AE2C431F3FDD4D
(IE4A74A61CDC56044C199B3C3D606B08E ), .I1CF1EE9FA60C0CDB15DD404CC8A269E5 (ICE73FC6522779AED50B02BB41E81D717 ), .I34F020684BFF4B1EAA406E693751B71D
(I25D595F391F999FD69AB7E7B5B1FA99C ), .IFB94B817F0BC84EC0734110F6EDE475A (IAE37CBAA4815C82EA96E8FA0802F7443 ), .I512A575E055CF9235066DBE4051242CB
(I50BD52F5094656ECEC3714E0BAE6B0DA ), .I391BF6A9C9F2ABEEA227F0E1F3F50A4F (IC781EE34DC62D08174F1793A9E3131B5 ), .IF0D7F78B99E50997A728E3731A197225
(I7568F6D9A53738CCE095CE231BAB3F85 ), .I9606837003EFA36A64A97C352D3D89A3 (ID23C9147B8CA6684051791F38B473984 ), .I4C1994114E1C49B9376320858F4E71F9
(ID873CC05798FE57AF43DD3C4E138769B ), .I2CB8399B2A61CDA9DB269D3567018E65 (I70E83CF258ED794C3E9EDE1260BF5578 ), .I46C5269B9FB24EF04CE2CC341C288EC7
(I46C5269B9FB24EF04CE2CC341C288EC7 ), .I3C9AD458B89B2FAABD743BF4E13BF421 (I3C9AD458B89B2FAABD743BF4E13BF421 ), .I73ABD5619A9FB885445AC1E288EAF7F8
(6), .IBDE0431C8F903800F409661F4F56FD80 (IB26EBF559CA483EACBAD1BCA4C580AF2 ) ) I79BD32F43383B22845A03B1C07DFF506
( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ),
.ICB680FEAB46B6D635CD9DD6BB49A6A20 (I8220BA29B6C07A3A107C2B3234F5FB06 ), .I8FF768DAF4C56D1B2D217B2C02B6D4EC (I7DA2457F5006629E45D78C4FC855DCF8 ),
.I9E5E6E86745F53F982BC3862031A206B (IBB764C0D62FD349F6FB3F52A8C78424E ), .I3AD72E1D6C16169DB8A27F1681293009 (IE074E5B8DF895724AB3B5023BAC298BC ),
.I0DE44F162EF92573C5DE1249527F6E9D (IDA2FA24095F53E4EBBAC1E30772082B4 ), .I2E9CC9AFC2E4742F852CB037CFC7E0A1 (I27FBA72EC841BBBDD25E028A08A3F06C ),
.I8B1798242C3B0E655181D0D365813614 (I8B1798242C3B0E655181D0D365813614 ), .IE145222FDBDC80109E12FA72D3D3C655 (IE145222FDBDC80109E12FA72D3D3C655 ),
.ID43AC1009727D128F1C5DFE4640CA5AB (ID43AC1009727D128F1C5DFE4640CA5AB ), .IB610431939CB8180EAC2403672BAF58D (IB610431939CB8180EAC2403672BAF58D ),
.I3C7A9FA839F554D8898020C4831479E2 (IC7DB18773990D347CEF55E672D6B2C05 ), .I74A0936EE8FD1443A2C6745A4F3F6B5E (I39A06B46F4E1C11EE4BFB781E3B4F32A ),
.I369BA2FFB5D41DF25F9BC3AB126D6607 (I369BA2FFB5D41DF25F9BC3AB126D6607 ), .I1C0271AD5E8E9E9164909E468AD0B212 (ID54A2FD9EE0AEAC4E7AC2A4D30D28B9B ),
.I6EC1BE4B18EC6AA3D88A5D45B614565E (I6EC1BE4B18EC6AA3D88A5D45B614565E [6]), .I56148DDDF284443347FFCF4F9C3BE61A (I81BF37FCB51B492DCA857F28ABD8D76E [6]),
.I24C403550AE065D7D1B7266142886226 (I24C403550AE065D7D1B7266142886226 ), .I438B8BD876741F9B46EB770E92F808B7 (I438B8BD876741F9B46EB770E92F808B7 [11:0]),
.I5FE75BE614D4F52DB327549B36203350 (I74CF4D6FE5B30BB30E40AFCA2A08A220 [6]), .I3D6C771D05CA1A769E61302C086494B8 (I3D6C771D05CA1A769E61302C086494B8 ),
.I357B3043EDACE3EBECE8F54D79B9F90A (I357B3043EDACE3EBECE8F54D79B9F90A ), .I0AAD559CF33A5CBA597990658774FEB3 (I0AAD559CF33A5CBA597990658774FEB3 ),
.I923204A95D8CBB206587CF32BEDCF4EF (I923204A95D8CBB206587CF32BEDCF4EF ), .ICF9D8FD31DFC7D20DAF939C6D75F1518 (ICF9D8FD31DFC7D20DAF939C6D75F1518 [6]),
.IDF550B17734BF16B7E410B19BB31E276 (IB9FE9C794CFE66C9E361CA5E0C2E0ED0 ), .I8ED9B9C1D9F58C5D06A9443AD901E8C6 (I200264A7B4F7EBBCB0636F8B0C705433 ),
.IA976D63BEECA80DCE31365CF56EC0248 (I5FCD09AF69B4D4969F86A3686036D558 ), .I5E3CE5AF5C34D232BFB139B63D9912B4 (IECF63199E2CFF774FC2362604C428EEF ),
.IBEF3E5F9395E2C7822AE03D6461DEBBB (IABDBB85ACD3277D447B4FD8665EA150B ), .I7E6CFD6A7DCAB9CD2188D044C7D716A6 (IB77F87CED77CEC2F6256375F35443CD0 ),
.I3A34691662384260F0524DD7F650E75A (IAF3303768435E5C76A60A5987AF1CD0A ), .IC2F58AB5028C1D2C53C6EF47A4975D0A (I2130A737A8CF0DAA0688CD61C692C53A ),
.I112E0A79129A8BC6DD4C13647C31F8A0 (I009BA1F74DBCC8E4177F1254D60DCAE9 ), .IE4B6DD43E04940631EF58BA04EA58997 (IACF97B89AE62537A26788BDFCE846ED1 [6]),
.I3A095084CDFDFA56A0E67616A78D3B25 (I01D4C6B20466D26621C6DA5816817455 [6]), .I81CD7F184DF8D58A1F2324E975A6816C (I46A701488EBE724B47736C3C7A47A876 [6]),
.I83C4A4200EB2B3F6766D338284ECAAAF (IFE63F76C2A46B87271596BE8D0FFD21A [6]), .I42A419EB6EB8D11234AC3B2BCA0AE593 (I3710541DAEAC21250982ECECA6E16679 ),
.IA41AC3CC6BC050DDC172724AB311315B (IEF2F499EA80B8075F4C485F59E3AA64D ), .I31CF69FF368B36B4D6612DF16B3ABC6B (I21EE6CA5EBC86B66AC5EE8AF763FB838 [6]),
.IFE4A8CBA73734C6F0F0A078027E053D4 (I386D96EE2FCEC8374B24F3017B94BD4D ), .ID7A2A8B1E9D92B60194D5FAFAAB15208 (I11E1C086CA3C13B481A5977B8AD8694F ),
.IF274FAF97F5BACD693913BB418717A9D (I5C58E3085FDB240D9A5DD64A9CD3A30B ), .ID95C13E7EE1CFE6A8743FF9E62C25873 (IE0683883BF201CF74ADDEE61816AAD96 ),
.IC58E411F24D810EF60A7B8638ABCC0BB (IF4776D1E9086F7D152D43C91A22BC985 ), .I89CFFA73C7546481B72B0FB06D799AEE (I176659D1476D3660538A1C22EFD75A83 ),
.I270ED686C2EF2C1C8B5B55EC4A5AAE84 (ID0B88392A9310E618D259D3AE74555DF ), .ID5CCD4858CB5CC1B2EDEC682C7DE5AAD (I2467937CC723EBC133B60C885A06C7A8 ),
.I7D901091F9E0741061C75B54467D48A0 (I3FC95340E6F01F64D548828DC3B2A0FE ) ); else begin assign ICF9D8FD31DFC7D20DAF939C6D75F1518 [6]
= 1'b0; assign IACF97B89AE62537A26788BDFCE846ED1 [6] = 1'b0; assign I01D4C6B20466D26621C6DA5816817455 [6] = 1'b0;
assign I46A701488EBE724B47736C3C7A47A876 [6] = 1'b0; assign IFE63F76C2A46B87271596BE8D0FFD21A [6] = 1'b0; assign
I21EE6CA5EBC86B66AC5EE8AF763FB838 [6] = 1'b0; assign IB9FE9C794CFE66C9E361CA5E0C2E0ED0 = 1'b0; assign I200264A7B4F7EBBCB0636F8B0C705433
= 1'b0; assign I5FCD09AF69B4D4969F86A3686036D558 = 1'b0; assign IECF63199E2CFF774FC2362604C428EEF = 1'b0; assign
IABDBB85ACD3277D447B4FD8665EA150B = 1'b0; assign IB77F87CED77CEC2F6256375F35443CD0 = 1'b0; assign IAF3303768435E5C76A60A5987AF1CD0A
= 1'b0; assign I2130A737A8CF0DAA0688CD61C692C53A = 1'b0; assign I009BA1F74DBCC8E4177F1254D60DCAE9 = 3'b0; assign
I3710541DAEAC21250982ECECA6E16679 = 3'b0; assign IEF2F499EA80B8075F4C485F59E3AA64D = 3'b0; assign I386D96EE2FCEC8374B24F3017B94BD4D
= 32'b0; assign I11E1C086CA3C13B481A5977B8AD8694F = 1'b0; assign I5C58E3085FDB240D9A5DD64A9CD3A30B = 1'b0; assign
IE0683883BF201CF74ADDEE61816AAD96 = 1'b0; assign IF4776D1E9086F7D152D43C91A22BC985 = 11'b0; assign I176659D1476D3660538A1C22EFD75A83
= 1'b0; assign ID0B88392A9310E618D259D3AE74555DF = 1'b0; assign I2467937CC723EBC133B60C885A06C7A8 = 1'b0; assign
I3FC95340E6F01F64D548828DC3B2A0FE = 32'b0; end endgenerate  generate if (I25B649490B20A1FEC9A1AA60AB0C6D5E ) I2296FC491415818D18357D6C2D700C14
# ( .IFC1FF746397E6A576E9FEB281890A248 (IFB72ECF29D30B02049C030502F330CE7 ), .IAF1DF965ED0D670C125D16FDF91B875B
(I7E6B00724A48BA5DD1C5E397542EDDC2 ), .IB7B379BA36F36F0638F4F33C7598CC85 (I5C146FC803FDD1163A6BAEA53E6C5468 ), .ID9DCCEB6B5B42C479CB9D2B3C992035D
(IE3404D24C7B1FA263F2EACB5CC85BFF6 ), .I251C6E5612F7B344EC3156CB9A93BE5B (IB23260A86DA99A28163B5E233CA42605 ), .ID7A688D3DA9A2C539FE87FC8998248CB
(IEF68A43ED89112E53191106DBA0EF113 ), .I96DBC3D130FB2B57DFB76E3E87DF89D2 (I95CE19A3BB94C8A24A8E3F3482EF6425 ), .I87B53E44EDBDCDA1796FB105323D3B17
(I7A84A5F1499409083F731D2A584D2D42 ), .IF9554E0938E353BDC05ABE0C628E3BE9 (I76069160333C4C8E92944FC3A3827ED6 ), .I37C708634F442A3B0568DA0BB576511F
(I8EF5BB87B22B910665D13A80C6724D14 ), .I7B125DA60401B7C86EB027E9E9262847 (IFA5339CE0FEDFF3B45CF3C0167564EA1 ), .I8BEE88809FA5712893BC59FF0E17ADB2
(ID3A400426A266A6F4E75F7686B9028CD ), .I7DF5A90920A562D09AA22D2DFA657124 (I071A2CF414FF8A814D779E1F54247BF1 ), .I0243B4A4E84E0712929C806F438E6AA9
(I3F7B58F167F56FB985F8908CA1B7E3AE ), .I7050B96C0C45A812BBFC45C2A30F272C (I62A26688D23065F69E9B9D6339AA01A5 ), .IB7C70D5D7B0DDF146F4D402BEE6F6FA6
(IE4774E19FB83A84DBF540368C45EA3A3 ), .I1CBD8B214B4765FBC7FA828F0C62BC94 (I5ACFA0E62CCC520EE4DA1BA399F1B7E6 ), .I677BE3663880CBE6E5AE2C431F3FDD4D
(IF1CB2B99D8669C68B68BC468C83323DF ), .I1CF1EE9FA60C0CDB15DD404CC8A269E5 (I245B45EC852C565EDD1AAC06E80DABD2 ), .I34F020684BFF4B1EAA406E693751B71D
(I59DF7AA363A19A361E3A844AD6039C40 ), .IFB94B817F0BC84EC0734110F6EDE475A (IAF2433492FE33171692143422229D319 ), .I512A575E055CF9235066DBE4051242CB
(I721D73CBB11DB0EC9DF361993F6A92EA ), .I391BF6A9C9F2ABEEA227F0E1F3F50A4F (IE0DA0C810288CC00DF1F3AE622FFB08F ), .IF0D7F78B99E50997A728E3731A197225
(IEB4CAA0AE4F26FAC1DAA6B9884179DEA ), .I9606837003EFA36A64A97C352D3D89A3 (I070D33CDFCF15FB7B4DD88019C0E39E2 ), .I4C1994114E1C49B9376320858F4E71F9
(I8302D4B9F46621BBB824B1CC96E2E724 ), .I2CB8399B2A61CDA9DB269D3567018E65 (I26BFDE09E6F548FBAC63338567411C7E ), .I46C5269B9FB24EF04CE2CC341C288EC7
(I46C5269B9FB24EF04CE2CC341C288EC7 ), .I3C9AD458B89B2FAABD743BF4E13BF421 (I3C9AD458B89B2FAABD743BF4E13BF421 ), .I73ABD5619A9FB885445AC1E288EAF7F8
(7), .IBDE0431C8F903800F409661F4F56FD80 (IB26EBF559CA483EACBAD1BCA4C580AF2 ) ) I854293011C70645A5B39295028B2D50B
( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ),
.ICB680FEAB46B6D635CD9DD6BB49A6A20 (I4FB68E387DB515A46DAA2DABF6E0D1D8 ), .I8FF768DAF4C56D1B2D217B2C02B6D4EC (IBA4DC2E68E546946B55995DB900F74F7 ),
.I9E5E6E86745F53F982BC3862031A206B (I28A9F4DDE0D0FFADF8668EFA99C6DA03 ), .I3AD72E1D6C16169DB8A27F1681293009 (IE02A2D602D1C83798270DD49EF6A4D23 ),
.I0DE44F162EF92573C5DE1249527F6E9D (I4DBB86A2215D89E37CDE4EC7DC8435C5 ), .I2E9CC9AFC2E4742F852CB037CFC7E0A1 (I8DCB72E575B62CC266039827C0238E34 ),
.I8B1798242C3B0E655181D0D365813614 (I8B1798242C3B0E655181D0D365813614 ), .IE145222FDBDC80109E12FA72D3D3C655 (IE145222FDBDC80109E12FA72D3D3C655 ),
.ID43AC1009727D128F1C5DFE4640CA5AB (ID43AC1009727D128F1C5DFE4640CA5AB ), .IB610431939CB8180EAC2403672BAF58D (IB610431939CB8180EAC2403672BAF58D ),
.I3C7A9FA839F554D8898020C4831479E2 (IC7DB18773990D347CEF55E672D6B2C05 ), .I74A0936EE8FD1443A2C6745A4F3F6B5E (I39A06B46F4E1C11EE4BFB781E3B4F32A ),
.I369BA2FFB5D41DF25F9BC3AB126D6607 (I369BA2FFB5D41DF25F9BC3AB126D6607 ), .I1C0271AD5E8E9E9164909E468AD0B212 (IA5469486BB0530B9AA1B819A3C7A9583 ),
.I6EC1BE4B18EC6AA3D88A5D45B614565E (I6EC1BE4B18EC6AA3D88A5D45B614565E [7]), .I56148DDDF284443347FFCF4F9C3BE61A (I81BF37FCB51B492DCA857F28ABD8D76E [7]),
.I24C403550AE065D7D1B7266142886226 (I24C403550AE065D7D1B7266142886226 ), .I438B8BD876741F9B46EB770E92F808B7 (I438B8BD876741F9B46EB770E92F808B7 [11:0]),
.I5FE75BE614D4F52DB327549B36203350 (I74CF4D6FE5B30BB30E40AFCA2A08A220 [7]), .I3D6C771D05CA1A769E61302C086494B8 (I3D6C771D05CA1A769E61302C086494B8 ),
.I357B3043EDACE3EBECE8F54D79B9F90A (I357B3043EDACE3EBECE8F54D79B9F90A ), .I0AAD559CF33A5CBA597990658774FEB3 (I0AAD559CF33A5CBA597990658774FEB3 ),
.I923204A95D8CBB206587CF32BEDCF4EF (I923204A95D8CBB206587CF32BEDCF4EF ), .ICF9D8FD31DFC7D20DAF939C6D75F1518 (ICF9D8FD31DFC7D20DAF939C6D75F1518 [7]),
.IDF550B17734BF16B7E410B19BB31E276 (IDEEB7827D919A8134F28A8BCC126AD5D ), .I8ED9B9C1D9F58C5D06A9443AD901E8C6 (IA7846F08DDB80EC63AA4A9EC1770A3F0 ),
.IA976D63BEECA80DCE31365CF56EC0248 (I93A8E9B4C6DB1D603A05A9591C4339C9 ), .I5E3CE5AF5C34D232BFB139B63D9912B4 (I17CB952AA0F6F5C6792E1381BEB60CA3 ),
.IBEF3E5F9395E2C7822AE03D6461DEBBB (IEB1DC53BA14A2028F346A4C10651DA08 ), .I7E6CFD6A7DCAB9CD2188D044C7D716A6 (I7616B3B0828958A3CA36203B840CF4D6 ),
.I3A34691662384260F0524DD7F650E75A (I246B1D75EEA1239D65C20304AF791CB4 ), .IC2F58AB5028C1D2C53C6EF47A4975D0A (IBCEA86C0BDF1E124E6697E40D620DD0A ),
.I112E0A79129A8BC6DD4C13647C31F8A0 (I11D20DB2F186022215040429BE705A72 ), .IE4B6DD43E04940631EF58BA04EA58997 (IACF97B89AE62537A26788BDFCE846ED1 [7]),
.I3A095084CDFDFA56A0E67616A78D3B25 (I01D4C6B20466D26621C6DA5816817455 [7]), .I81CD7F184DF8D58A1F2324E975A6816C (I46A701488EBE724B47736C3C7A47A876 [7]),
.I83C4A4200EB2B3F6766D338284ECAAAF (IFE63F76C2A46B87271596BE8D0FFD21A [7]), .I42A419EB6EB8D11234AC3B2BCA0AE593 (I73B39CB9A73EAB03AD04B21F62F95224 ),
.IA41AC3CC6BC050DDC172724AB311315B (I700C2FF696E95E1F0C6E6B8EB54971BC ), .I31CF69FF368B36B4D6612DF16B3ABC6B (I21EE6CA5EBC86B66AC5EE8AF763FB838 [7]),
.IFE4A8CBA73734C6F0F0A078027E053D4 (I49850943EA73C8BE46401A2FC9B67D74 ), .ID7A2A8B1E9D92B60194D5FAFAAB15208 (I14F6DF0BCAC12F6EBAD7145BDD4B2D26 ),
.IF274FAF97F5BACD693913BB418717A9D (IB85FB30E34AF0B105FD21BBBB73605EA ), .ID95C13E7EE1CFE6A8743FF9E62C25873 (IE67F175E6F2CC66DDCAD62CCD21F3551 ),
.IC58E411F24D810EF60A7B8638ABCC0BB (I58A4869C5AA5FC57B207E7883C179856 ), .I89CFFA73C7546481B72B0FB06D799AEE (I9DD533FE3D53A79078BF27CC1058785B ),
.I270ED686C2EF2C1C8B5B55EC4A5AAE84 (I4D0BD33FE293DDEE3A568B64EE8F63F1 ), .ID5CCD4858CB5CC1B2EDEC682C7DE5AAD (I42FFAA9F6065323EF66FBE15FAE57258 ),
.I7D901091F9E0741061C75B54467D48A0 (IE8EF8CF3D14B7C15DC96E6E2DC4BA14A ) ); else begin assign ICF9D8FD31DFC7D20DAF939C6D75F1518 [7]
= 1'b0; assign IACF97B89AE62537A26788BDFCE846ED1 [7] = 1'b0; assign I01D4C6B20466D26621C6DA5816817455 [7] = 1'b0;
assign I46A701488EBE724B47736C3C7A47A876 [7] = 1'b0; assign IFE63F76C2A46B87271596BE8D0FFD21A [7] = 1'b0; assign
I21EE6CA5EBC86B66AC5EE8AF763FB838 [7] = 1'b0; assign IDEEB7827D919A8134F28A8BCC126AD5D = 1'b0; assign IA7846F08DDB80EC63AA4A9EC1770A3F0
= 1'b0; assign I93A8E9B4C6DB1D603A05A9591C4339C9 = 1'b0; assign I17CB952AA0F6F5C6792E1381BEB60CA3 = 1'b0; assign
IEB1DC53BA14A2028F346A4C10651DA08 = 1'b0; assign I7616B3B0828958A3CA36203B840CF4D6 = 1'b0; assign I246B1D75EEA1239D65C20304AF791CB4
= 1'b0; assign IBCEA86C0BDF1E124E6697E40D620DD0A = 1'b0; assign I11D20DB2F186022215040429BE705A72 = 3'b0; assign
I73B39CB9A73EAB03AD04B21F62F95224 = 3'b0; assign I700C2FF696E95E1F0C6E6B8EB54971BC = 3'b0; assign I49850943EA73C8BE46401A2FC9B67D74
= 32'b0; assign I14F6DF0BCAC12F6EBAD7145BDD4B2D26 = 1'b0; assign IB85FB30E34AF0B105FD21BBBB73605EA = 1'b0; assign
IE67F175E6F2CC66DDCAD62CCD21F3551 = 1'b0; assign I58A4869C5AA5FC57B207E7883C179856 = 11'b0; assign I9DD533FE3D53A79078BF27CC1058785B
= 1'b0; assign I4D0BD33FE293DDEE3A568B64EE8F63F1 = 1'b0; assign I42FFAA9F6065323EF66FBE15FAE57258 = 1'b0; assign
IE8EF8CF3D14B7C15DC96E6E2DC4BA14A = 32'b0; end endgenerate  IF8888DF840520FCED3157D151D128B3B #( .IE50492CEE03959C13AD5E521CC7F2FEF
(IE50492CEE03959C13AD5E521CC7F2FEF ), .I0B3C14F69FAC563649E26679A3D8B1CD (I0B3C14F69FAC563649E26679A3D8B1CD ), .IFA272F301A5935EE15CB134524665363
(IFA272F301A5935EE15CB134524665363 ), .IE690B7723F136DA02896C0728DDADB49 (IE690B7723F136DA02896C0728DDADB49 ), .I55BE27080C370AF723A4FE096014E875
(I55BE27080C370AF723A4FE096014E875 ), .IB2560D175E4507798B84D6E659FD6373 (IB2560D175E4507798B84D6E659FD6373 ), .I25B649490B20A1FEC9A1AA60AB0C6D5E
(I25B649490B20A1FEC9A1AA60AB0C6D5E ) ) I4108110328C413276966776688BEAB97 ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ),
.I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .IE145222FDBDC80109E12FA72D3D3C655 (IE145222FDBDC80109E12FA72D3D3C655 ),
.I2AD6292CA4A68298ECB0EB04E60DC338 (I60003168A46706B958CCEC72E50AC23E ), .I7E1B3386EACDCC0730096B4BEBD3FC11 (I111827C337F00C09A8C61C3DCE514338 ),
.IE10AAAB7732A262D17819D08F8A724BC (ICF847A44ADAE70C9998962202A23AB4E ), .IDF7BAD8C79D202960378A7387FEE4794 (IC4C35B8C650EEF422BEF8C68B5A9359D ),
.I57990336F36AA63E9FBA5533A4E25FA3 (IB624795CEFFC2094E111CAD5578DAE1C ), .IED35F37F7AD8CD8C1B242C9C79E11FA3 (IB56580C539321C40E6B44EB394A9EECF ),
.ID2BF5B6DEE97B309004C8AC7C3F5B8B3 (I400149787F2546E3D0331041FB8123FC ), .I3C7A9FA839F554D8898020C4831479E2 (I3C7A9FA839F554D8898020C4831479E2 ),
.I74A0936EE8FD1443A2C6745A4F3F6B5E (I74A0936EE8FD1443A2C6745A4F3F6B5E ), .I369BA2FFB5D41DF25F9BC3AB126D6607 (I369BA2FFB5D41DF25F9BC3AB126D6607 ),
.I2CB69D0EFAF8ADA6B6211F64BA9D2B52 (IACF97B89AE62537A26788BDFCE846ED1 ), .I3EEF1AC61F6E4A2B704EBA11EF949965 (I01D4C6B20466D26621C6DA5816817455 ),
.I25EC384599199AF35E4D0B3B873187EF (I46A701488EBE724B47736C3C7A47A876 ), .I8F57B8D98905C89F4D3B91CA626C25BA (IFE63F76C2A46B87271596BE8D0FFD21A ),
.I56148DDDF284443347FFCF4F9C3BE61A (I81BF37FCB51B492DCA857F28ABD8D76E [8]), .I24C403550AE065D7D1B7266142886226 (I24C403550AE065D7D1B7266142886226 ),
.I5FE75BE614D4F52DB327549B36203350 (I5FE75BE614D4F52DB327549B36203350 ), .I0AAD559CF33A5CBA597990658774FEB3 (I0AAD559CF33A5CBA597990658774FEB3 ),
.I923204A95D8CBB206587CF32BEDCF4EF (I923204A95D8CBB206587CF32BEDCF4EF ), .I20CD33DEFBDF51E2A5352736B083738D (I20CD33DEFBDF51E2A5352736B083738D ),
.I8ED9B9C1D9F58C5D06A9443AD901E8C6 (I18AB4B503F92B00D610DFDE3078A4B8F ), .IA976D63BEECA80DCE31365CF56EC0248 (IAF7DC8691D3941B7E52C532F1E8C7FE1 ),
.I5E3CE5AF5C34D232BFB139B63D9912B4 (IBFA78112A3EFE7AB665D3E3A9A588B1D ), .IBEF3E5F9395E2C7822AE03D6461DEBBB (I94288AE7E6EFEA1989E284E9B2867097 ),
.I7E6CFD6A7DCAB9CD2188D044C7D716A6 (IDEB44FD98C3E74E285A47A4BD69A7619 ), .I3A34691662384260F0524DD7F650E75A (I3A3A0FDF754EB1C6D50FABC25DBFC696 ),
.IC2F58AB5028C1D2C53C6EF47A4975D0A (ICCD7B28178C3803739C5C1C758B836E2 ), .ID3E7F4B58943229FEE6313A36B3F8693 (IC7DB18773990D347CEF55E672D6B2C05 ),
.I1FDEC1735547330C00A0B8DFE1FB10C3 (I39A06B46F4E1C11EE4BFB781E3B4F32A ), .I439AF6D496491F5F7C23217209B43C31 (IA513FFA7CDD6BF8E65B629CB494239A4 ),
.IFE4A8CBA73734C6F0F0A078027E053D4 (I6DFBACFF2E5A466B93A00001848429F7 ), .ID7A2A8B1E9D92B60194D5FAFAAB15208 (I7CA41EFBA3D0548B989711570EA40B95 ),
.IF274FAF97F5BACD693913BB418717A9D (IC30C68A9857DD63CE5A51E5943CEB3AF ), .ID95C13E7EE1CFE6A8743FF9E62C25873 (I8824AFA21C1B61513D8DE94591B948FB ),
.I0DA874BD2204FA5231F61AC696D6584A (IB5292E1DAB3B0E7E62E43F792E80D8F1 ), .I270ED686C2EF2C1C8B5B55EC4A5AAE84 (ID4282AD4BEFA96986B17E55149DF417C )
);  IFF5E0986AB6F727F3EEDED75702CE45A # ( .IAB32DAC10CBDBE04FD5EDBF7A576CAF9 (IAB32DAC10CBDBE04FD5EDBF7A576CAF9 ),
.I5F8A137EF3A5FDA6F2493F06E8FA441C (IE3D0FF95EEFE7CF51F7D6968D26EAB4A ), .I66C185998F46A7148163982E39BCD296 (I66C185998F46A7148163982E39BCD296 )
) IE0EBA42E51B882F4CBD779D6D5FBF73E ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .I3FF97406B3ED373B267711109A980AF9 (I3FF97406B3ED373B267711109A980AF9 ), .I91C25096707DEBEF0FC17788A26B01A1
(I56519DD369C66F1A0EA1EE3D2398E0EF ), .I6777AFB972CFFDA974EE962374CC84A0 (IC0667A37FE3E5F8D3579C6AEF86F5C24 ), .IA29FAC409EB1AFED4EA6D47BD6948E58
(IB907C2624CE144BCE5A772623C46F678 ), .I39B913343A3C8C7ED94053B14CAC4B0B ( ), .ID721B306FF47217933BAF6C84043D7D0
(I81BF37FCB51B492DCA857F28ABD8D76E ) ); endmodule 
 `timescale 1 ns / 1 ps
module IA8C351750B9DBEE4D8ADA94748C8E5D1 # (parameter I61D0345D311EC6FFC08DDDECE5F6127A = 256, parameter I5C6C6CD7723900C21B3A76E887CEE164
= 32, parameter I64BB723AC8F87F7AEBA73BF190ED5F8F = 32 ) ( input wire ICCFB0F435B37370076102F325BC08D20 , input
wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire I8F36BEAA79ADAC31FBCBAC1B805C772E , input wire IE52544EAEF6757A8A982FC14CE507F8C ,
input wire [9:0] IAC8BFFA8C250FC35278EA36BA7C00B42 , input wire [1:0] I27CF4DD7FCBC7E0A229344EDF94F2651 , input
wire I1A55EB74BDB9184AA980B07905C85479 , input wire IC79EC9A9F373F4B71374BDF6EDD31DE6 , input wire ID8853B025150C80EE45BBA98E5BEA3A8 ,
input wire [I5C6C6CD7723900C21B3A76E887CEE164 - 1:0] I04BC24D2B6403E54A64DE9E6C9ABAA2B , input wire I3F6FB755DC9826D564C143FF9E32F032 ,
input wire IE315CDCA06C9620D5C0AB966E553F0C3 , output wire [$clog2(I61D0345D311EC6FFC08DDDECE5F6127A ) - 1:0] I7740E93179670969593F64CBA98864D9 ,
output wire [$clog2(I61D0345D311EC6FFC08DDDECE5F6127A ) - 1:0] I89011D8BA1FC92A73CD875E098FE685C , output wire [I64BB723AC8F87F7AEBA73BF190ED5F8F :0]
I7D649F765882BD862315E777ABA5263F , output wire I87AD4A36141619A102AD5166323D80AB , output wire [$clog2(I61D0345D311EC6FFC08DDDECE5F6127A
+ 1) - 1:0] ID7FCE45A65ADDB17F91F73A1B506BB5B , output wire I8BB939FF2AFDE7B2A1E480DCB61CE354 , output wire I585F74DE05DD9C1C7070D6B4F6E181C2 ,
output wire [$clog2((I61D0345D311EC6FFC08DDDECE5F6127A * (I64BB723AC8F87F7AEBA73BF190ED5F8F /I5C6C6CD7723900C21B3A76E887CEE164 ))
+ 1) - 1:0] I233E0C0C8E5150F0CD8258F276D93942 , output wire IBE0D6810EBD63B5C428623C578CF6D3A );  localparam IFA55551D85BC21F7BB69A4B7EF5E7D87
= I64BB723AC8F87F7AEBA73BF190ED5F8F / I5C6C6CD7723900C21B3A76E887CEE164 ; localparam IC95B888EAB7163F28FD516505CC99B4A
= 2'b00; localparam I33391FACE7091AC60C06B63939F2297C = 2'b01; localparam IB2A3AE77A1D62E86F85DC16314DCC934 = 2'b10;
localparam IA05DD9BECCC202CEB5D936A7AE596D73 = 2'b11; localparam I823055679D0D42FB8C0624248C03ECD8 = $clog2(I61D0345D311EC6FFC08DDDECE5F6127A );
localparam IC17027476895C8A3932B682A6B268544 = (IFA55551D85BC21F7BB69A4B7EF5E7D87 == 1) ? ($clog2(IFA55551D85BC21F7BB69A4B7EF5E7D87 )
+ 1) : $clog2(IFA55551D85BC21F7BB69A4B7EF5E7D87 ); localparam I05264B2FA834FBEA729752C27B778963 = $clog2(I61D0345D311EC6FFC08DDDECE5F6127A
+ 1); localparam I6BAD12625217B36EDD0324B5AD4BB875 = $clog2((I61D0345D311EC6FFC08DDDECE5F6127A * IFA55551D85BC21F7BB69A4B7EF5E7D87 )
+ 1);  reg [IC17027476895C8A3932B682A6B268544 - 1:0] I10F60E589450CD09FF7A498641DE26F8 ; reg IDA82F4C78A43B62E1C09ED19A1443221 ;
reg IF4B2F356412545C21578876129150C2F ; reg [10:0] I86FE3F5063E3F8D29DC1B4511B190C1F ; reg I1894079D486CFFF5D3FD4A0BD4CF0823 ;
reg I149E6E0597FD4E21363A409D472C2961 ; reg [I823055679D0D42FB8C0624248C03ECD8 - 1:0] I3283453B42BD77672B8ACE724ACDA314 ;
reg I7443F8A38FD149075A7DFFAF8C0D2BE9 ; reg [I823055679D0D42FB8C0624248C03ECD8 - 1:0] IF8FA22381AE98928C01C1A8EF2CB0DC6 ;
reg [I64BB723AC8F87F7AEBA73BF190ED5F8F - 1:0] I690EDD8A1FA9E66FB9012E57D65F740E ; reg I68525D8B661ABC93EC5BB1B92FE9724E ;
reg IC884C37BE792A5FAFAED7FC0B3F66BCD ; reg [10:0] I1A31CF65341BC1BA21B167CA7607B766 ; reg [1:0] I3C78D9AB59D6164851A819C5BA6C7C04 ;
reg [2:0] IC62A92297514890D9C19621875B887EF ; reg I49AAD9C7D99712758382319F50D699DA ; reg IE31D0AF3EFB3124913CD965CEE542B24 ;
reg [I05264B2FA834FBEA729752C27B778963 - 1:0] IDDFF27981262750D43304A01A2EBF659 ; reg I05305DB38B053FE192F0B71598347D85 ;
reg [I6BAD12625217B36EDD0324B5AD4BB875 - 1:0] IE1A203A1BCBBA5F947F638C3DFB65BF8 ; wire I2C3263714ADF8DC5044612F1D1CA7C60 ;
wire [I64BB723AC8F87F7AEBA73BF190ED5F8F :0] I37967D3D367DBC529BC9A9CCD8D412C3 ; wire IB571869C20EDD4E0FBF88724DD731261 ;
wire [I64BB723AC8F87F7AEBA73BF190ED5F8F - 1:0] I8AC98A8524CB0CAD513AB7EAD12AB430 ; wire I82A06AFC4695660C2A666925552E8623 ;
wire [10:0] I181D2D586A16E282B74A78EECE6F0DFB ; wire IFBDC6122402AF53F2C50F690FE464A6B ; wire I8CAAE4487A3778130CA1C80C5F36EE61 ;
 assign I7740E93179670969593F64CBA98864D9 = I3283453B42BD77672B8ACE724ACDA314 ; assign I89011D8BA1FC92A73CD875E098FE685C
= IF8FA22381AE98928C01C1A8EF2CB0DC6 ; assign I7D649F765882BD862315E777ABA5263F = (I5C6C6CD7723900C21B3A76E887CEE164
== I64BB723AC8F87F7AEBA73BF190ED5F8F ) ? {I3F6FB755DC9826D564C143FF9E32F032 , I04BC24D2B6403E54A64DE9E6C9ABAA2B }
: I37967D3D367DBC529BC9A9CCD8D412C3 ; assign I87AD4A36141619A102AD5166323D80AB = IB571869C20EDD4E0FBF88724DD731261 ;
assign ID7FCE45A65ADDB17F91F73A1B506BB5B = IDDFF27981262750D43304A01A2EBF659 ; assign I8BB939FF2AFDE7B2A1E480DCB61CE354
= I1894079D486CFFF5D3FD4A0BD4CF0823 ; assign I585F74DE05DD9C1C7070D6B4F6E181C2 = I05305DB38B053FE192F0B71598347D85 ;
assign I233E0C0C8E5150F0CD8258F276D93942 = IE1A203A1BCBBA5F947F638C3DFB65BF8 ; assign IBE0D6810EBD63B5C428623C578CF6D3A
= I149E6E0597FD4E21363A409D472C2961 ;  assign I2C3263714ADF8DC5044612F1D1CA7C60 = (ID8853B025150C80EE45BBA98E5BEA3A8
| IFBDC6122402AF53F2C50F690FE464A6B ) & !I1894079D486CFFF5D3FD4A0BD4CF0823 ; assign IB571869C20EDD4E0FBF88724DD731261
= (I5C6C6CD7723900C21B3A76E887CEE164 == I64BB723AC8F87F7AEBA73BF190ED5F8F ) ? I8CAAE4487A3778130CA1C80C5F36EE61
: I82A06AFC4695660C2A666925552E8623 ; assign I82A06AFC4695660C2A666925552E8623 = (I10F60E589450CD09FF7A498641DE26F8
== (IFA55551D85BC21F7BB69A4B7EF5E7D87 - 1)) ? I8CAAE4487A3778130CA1C80C5F36EE61 : (I8CAAE4487A3778130CA1C80C5F36EE61
& I3F6FB755DC9826D564C143FF9E32F032 ); assign I181D2D586A16E282B74A78EECE6F0DFB = (IDA82F4C78A43B62E1C09ED19A1443221 )
? ((IF4B2F356412545C21578876129150C2F ) ? I86FE3F5063E3F8D29DC1B4511B190C1F + 4 : I86FE3F5063E3F8D29DC1B4511B190C1F
+ 3) : ((IF4B2F356412545C21578876129150C2F ) ? {11{1'b0}} + 4 : {11{1'b0}} + 3); assign IFBDC6122402AF53F2C50F690FE464A6B
= (I1A55EB74BDB9184AA980B07905C85479 & ~I49AAD9C7D99712758382319F50D699DA & ~I1894079D486CFFF5D3FD4A0BD4CF0823 )
| (I49AAD9C7D99712758382319F50D699DA & IE31D0AF3EFB3124913CD965CEE542B24 & ~I1894079D486CFFF5D3FD4A0BD4CF0823 );
assign I8CAAE4487A3778130CA1C80C5F36EE61 = IE315CDCA06C9620D5C0AB966E553F0C3 & !I149E6E0597FD4E21363A409D472C2961 ;
 generate if (IFA55551D85BC21F7BB69A4B7EF5E7D87 == 1) begin assign I37967D3D367DBC529BC9A9CCD8D412C3 = {I3F6FB755DC9826D564C143FF9E32F032 ,
I04BC24D2B6403E54A64DE9E6C9ABAA2B }; end endgenerate generate if (IFA55551D85BC21F7BB69A4B7EF5E7D87 == 2) begin
assign I37967D3D367DBC529BC9A9CCD8D412C3 = {I3F6FB755DC9826D564C143FF9E32F032 , ((I3F6FB755DC9826D564C143FF9E32F032
&& (I10F60E589450CD09FF7A498641DE26F8 == 0)) ? I04BC24D2B6403E54A64DE9E6C9ABAA2B : I690EDD8A1FA9E66FB9012E57D65F740E [I5C6C6CD7723900C21B3A76E887CEE164
- 1:0]), I04BC24D2B6403E54A64DE9E6C9ABAA2B }; end endgenerate generate if (I64BB723AC8F87F7AEBA73BF190ED5F8F > I5C6C6CD7723900C21B3A76E887CEE164 )
assign I8AC98A8524CB0CAD513AB7EAD12AB430 = {I690EDD8A1FA9E66FB9012E57D65F740E [I64BB723AC8F87F7AEBA73BF190ED5F8F
- I5C6C6CD7723900C21B3A76E887CEE164 - 1:0], I04BC24D2B6403E54A64DE9E6C9ABAA2B }; else assign I8AC98A8524CB0CAD513AB7EAD12AB430
= I04BC24D2B6403E54A64DE9E6C9ABAA2B ; endgenerate  generate if (1'b1) begin : I8CDDE92DE2910086C77F2B20C50D61C7
reg [1:0] I102EDFAABB65014FC78C55AF4345F765 ; reg [1:0] ICA80E74165E79AFA565A1A052BE49F09 ; task I8BE101CBEF6D2810BAC0C6F6AC8DA3B8 ;
begin I10F60E589450CD09FF7A498641DE26F8 <= {IC17027476895C8A3932B682A6B268544 {1'b0}}; I1894079D486CFFF5D3FD4A0BD4CF0823
<= 1'b1; I149E6E0597FD4E21363A409D472C2961 <= 1'b0; I3283453B42BD77672B8ACE724ACDA314 <= 0; I7443F8A38FD149075A7DFFAF8C0D2BE9
<= 1'b0; IF8FA22381AE98928C01C1A8EF2CB0DC6 <= 0; IDDFF27981262750D43304A01A2EBF659 <= 0; IE1A203A1BCBBA5F947F638C3DFB65BF8
<= I61D0345D311EC6FFC08DDDECE5F6127A * IFA55551D85BC21F7BB69A4B7EF5E7D87 ; end endtask always @(posedge ICCFB0F435B37370076102F325BC08D20
or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin if (I9ED2A9117D3AEAF54CBA7AD69083BCB7 == 1'b0) begin I8BE101CBEF6D2810BAC0C6F6AC8DA3B8 ;
IDA82F4C78A43B62E1C09ED19A1443221 <= 1'b0; IF4B2F356412545C21578876129150C2F <= 1'b0; I86FE3F5063E3F8D29DC1B4511B190C1F
<= {11{1'b0}}; I690EDD8A1FA9E66FB9012E57D65F740E <= {I64BB723AC8F87F7AEBA73BF190ED5F8F {1'b0}}; I68525D8B661ABC93EC5BB1B92FE9724E
<= 1'b0; IC884C37BE792A5FAFAED7FC0B3F66BCD <= 1'b0; I3C78D9AB59D6164851A819C5BA6C7C04 <= 2'b0; IC62A92297514890D9C19621875B887EF
<= 3'b0; I49AAD9C7D99712758382319F50D699DA <= 1'b0; IE31D0AF3EFB3124913CD965CEE542B24 <= 1'b0; I05305DB38B053FE192F0B71598347D85
<= 1'b0; end else begin IDA82F4C78A43B62E1C09ED19A1443221 <= IE52544EAEF6757A8A982FC14CE507F8C ; IF4B2F356412545C21578876129150C2F
<= I8F36BEAA79ADAC31FBCBAC1B805C772E ; I86FE3F5063E3F8D29DC1B4511B190C1F <= {~(|IAC8BFFA8C250FC35278EA36BA7C00B42 ),
IAC8BFFA8C250FC35278EA36BA7C00B42 }; I3C78D9AB59D6164851A819C5BA6C7C04 <= I27CF4DD7FCBC7E0A229344EDF94F2651 ; if
(I1A55EB74BDB9184AA980B07905C85479 | I49AAD9C7D99712758382319F50D699DA ) begin if (IFBDC6122402AF53F2C50F690FE464A6B )
if (I1A31CF65341BC1BA21B167CA7607B766 > 2) I1A31CF65341BC1BA21B167CA7607B766 <= I1A31CF65341BC1BA21B167CA7607B766
- IFA55551D85BC21F7BB69A4B7EF5E7D87 ; else I1A31CF65341BC1BA21B167CA7607B766 <= {11{1'b0}}; end else I1A31CF65341BC1BA21B167CA7607B766
<= I181D2D586A16E282B74A78EECE6F0DFB ; if (IC79EC9A9F373F4B71374BDF6EDD31DE6 == 1'b1) I8BE101CBEF6D2810BAC0C6F6AC8DA3B8 ;
else begin if (I1A55EB74BDB9184AA980B07905C85479 | IE31D0AF3EFB3124913CD965CEE542B24 ) begin IE31D0AF3EFB3124913CD965CEE542B24
<= (I3C78D9AB59D6164851A819C5BA6C7C04 == IC95B888EAB7163F28FD516505CC99B4A ) ? 1'b1 : 1'b0; case (I3C78D9AB59D6164851A819C5BA6C7C04 )
I33391FACE7091AC60C06B63939F2297C : begin IC62A92297514890D9C19621875B887EF <= 3'b001; end IB2A3AE77A1D62E86F85DC16314DCC934
: begin IC62A92297514890D9C19621875B887EF <= 3'b011; end IA05DD9BECCC202CEB5D936A7AE596D73 : begin IC62A92297514890D9C19621875B887EF
<= 3'b111; end default : begin IC62A92297514890D9C19621875B887EF <= 3'b000; end endcase end else begin IC62A92297514890D9C19621875B887EF
<= (I3C78D9AB59D6164851A819C5BA6C7C04 == IC95B888EAB7163F28FD516505CC99B4A ) ? 3'b000 : (IC62A92297514890D9C19621875B887EF
- 1); IE31D0AF3EFB3124913CD965CEE542B24 <= (I3C78D9AB59D6164851A819C5BA6C7C04 == IC95B888EAB7163F28FD516505CC99B4A )
? 1'b1 : ((IC62A92297514890D9C19621875B887EF == 3'b001) ? 1'b1 : 1'b0); end  if (I8CAAE4487A3778130CA1C80C5F36EE61 )
begin I10F60E589450CD09FF7A498641DE26F8 <= ((I10F60E589450CD09FF7A498641DE26F8 == (IFA55551D85BC21F7BB69A4B7EF5E7D87
- 1)) || I3F6FB755DC9826D564C143FF9E32F032 ) ? {IC17027476895C8A3932B682A6B268544 {1'b0}} : (I10F60E589450CD09FF7A498641DE26F8
+ 1); I690EDD8A1FA9E66FB9012E57D65F740E <= I8AC98A8524CB0CAD513AB7EAD12AB430 ; end  I102EDFAABB65014FC78C55AF4345F765
= {I2C3263714ADF8DC5044612F1D1CA7C60 , IB571869C20EDD4E0FBF88724DD731261 }; case (I102EDFAABB65014FC78C55AF4345F765 )
2'b01: begin I1894079D486CFFF5D3FD4A0BD4CF0823 <= 1'b0; I7443F8A38FD149075A7DFFAF8C0D2BE9 <= I1894079D486CFFF5D3FD4A0BD4CF0823 ;
IDDFF27981262750D43304A01A2EBF659 <= IDDFF27981262750D43304A01A2EBF659 + 1; end 2'b10: begin I1894079D486CFFF5D3FD4A0BD4CF0823
<= I1894079D486CFFF5D3FD4A0BD4CF0823 | ((IDDFF27981262750D43304A01A2EBF659 == 1) ? 1'b1 : 1'b0); I7443F8A38FD149075A7DFFAF8C0D2BE9
<= (IDDFF27981262750D43304A01A2EBF659 == 2) ? 1'b1 : 1'b0; IDDFF27981262750D43304A01A2EBF659 <= IDDFF27981262750D43304A01A2EBF659
- 1; end endcase  ICA80E74165E79AFA565A1A052BE49F09 = {I2C3263714ADF8DC5044612F1D1CA7C60 , IB571869C20EDD4E0FBF88724DD731261 };
case (ICA80E74165E79AFA565A1A052BE49F09 ) 2'b01: begin I149E6E0597FD4E21363A409D472C2961 <= I149E6E0597FD4E21363A409D472C2961
| ((IE1A203A1BCBBA5F947F638C3DFB65BF8 == 1) ? 1'b1 : 1'b0); IE1A203A1BCBBA5F947F638C3DFB65BF8 <= IE1A203A1BCBBA5F947F638C3DFB65BF8
- IFA55551D85BC21F7BB69A4B7EF5E7D87 ; end 2'b10: begin I149E6E0597FD4E21363A409D472C2961 <= 1'b0; IE1A203A1BCBBA5F947F638C3DFB65BF8
<= IE1A203A1BCBBA5F947F638C3DFB65BF8 + IFA55551D85BC21F7BB69A4B7EF5E7D87 ; end endcase  I68525D8B661ABC93EC5BB1B92FE9724E
<= I2C3263714ADF8DC5044612F1D1CA7C60 ; IC884C37BE792A5FAFAED7FC0B3F66BCD <= (~I1894079D486CFFF5D3FD4A0BD4CF0823
& ~I2C3263714ADF8DC5044612F1D1CA7C60 ) | (IC884C37BE792A5FAFAED7FC0B3F66BCD & ~I68525D8B661ABC93EC5BB1B92FE9724E )
| (I68525D8B661ABC93EC5BB1B92FE9724E & ~I1894079D486CFFF5D3FD4A0BD4CF0823 ); I49AAD9C7D99712758382319F50D699DA <=
(I1A55EB74BDB9184AA980B07905C85479 & ~I49AAD9C7D99712758382319F50D699DA ) | (I49AAD9C7D99712758382319F50D699DA &
((I1A31CF65341BC1BA21B167CA7607B766 > IFA55551D85BC21F7BB69A4B7EF5E7D87 ) ? 1'b1 : ~IE31D0AF3EFB3124913CD965CEE542B24 ));
I05305DB38B053FE192F0B71598347D85 <= I68525D8B661ABC93EC5BB1B92FE9724E & IC884C37BE792A5FAFAED7FC0B3F66BCD ; if
(I2C3263714ADF8DC5044612F1D1CA7C60 == 1'b1) I3283453B42BD77672B8ACE724ACDA314 <= I3283453B42BD77672B8ACE724ACDA314
+ 1; if (IB571869C20EDD4E0FBF88724DD731261 == 1'b1) IF8FA22381AE98928C01C1A8EF2CB0DC6 <= IF8FA22381AE98928C01C1A8EF2CB0DC6
+ 1; end  end  end  end  endgenerate endmodule 
  `timescale 1 ns / 1 ps 
module I6433000F3EF06E04177C32D16C534889 # (parameter IB71844FFA3AB85FEF45EAB4D35395752 = 512, parameter I5C6C6CD7723900C21B3A76E887CEE164
= 32, parameter I64BB723AC8F87F7AEBA73BF190ED5F8F = 32, parameter I66C185998F46A7148163982E39BCD296 = "ecp3" ) (
input wire ICCFB0F435B37370076102F325BC08D20 , input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire [1:0] I27CF4DD7FCBC7E0A229344EDF94F2651 ,
input wire I1A55EB74BDB9184AA980B07905C85479 , input wire I48D61F5A0B5732A58912433B42CD9D0C , input wire [I5C6C6CD7723900C21B3A76E887CEE164
- 1:0] I04BC24D2B6403E54A64DE9E6C9ABAA2B , input wire I3F6FB755DC9826D564C143FF9E32F032 , input wire IE315CDCA06C9620D5C0AB966E553F0C3 ,
output wire [$clog2(IB71844FFA3AB85FEF45EAB4D35395752 + 1) - 1:0] ID7FCE45A65ADDB17F91F73A1B506BB5B , output wire
[I64BB723AC8F87F7AEBA73BF190ED5F8F - 1:0] I125028C7446331521D0434C10E8B0007 , output wire I8BB939FF2AFDE7B2A1E480DCB61CE354 ,
output wire IC9DE8233C6B1ADF4418EEF5B1F14BE49 , output wire I585F74DE05DD9C1C7070D6B4F6E181C2 , output wire [$clog2((IB71844FFA3AB85FEF45EAB4D35395752
* (I64BB723AC8F87F7AEBA73BF190ED5F8F /I5C6C6CD7723900C21B3A76E887CEE164 )) + 1) - 1:0] I233E0C0C8E5150F0CD8258F276D93942 ,
output wire IBE0D6810EBD63B5C428623C578CF6D3A );  localparam integer I36A1B4EB5B5564A6ED7EA4D42856EFB4 = $clog2(IB71844FFA3AB85FEF45EAB4D35395752 );
localparam integer I05264B2FA834FBEA729752C27B778963 = $clog2(IB71844FFA3AB85FEF45EAB4D35395752 + 1); localparam
integer I6BAD12625217B36EDD0324B5AD4BB875 = $clog2((IB71844FFA3AB85FEF45EAB4D35395752 * (I64BB723AC8F87F7AEBA73BF190ED5F8F /I5C6C6CD7723900C21B3A76E887CEE164 ))
+ 1); localparam integer IEC3803494FB0D58F44099BF28643CCC0 = I5C6C6CD7723900C21B3A76E887CEE164 + 1; localparam integer
I05F95435FA8D508B4820D9E064382614 = I64BB723AC8F87F7AEBA73BF190ED5F8F + 1; localparam integer IFA55551D85BC21F7BB69A4B7EF5E7D87
= I64BB723AC8F87F7AEBA73BF190ED5F8F / I5C6C6CD7723900C21B3A76E887CEE164 ;  wire [I05F95435FA8D508B4820D9E064382614
- 1:0] IFAF7F03355554E59A3861F8A72D71CA5 ; wire [I36A1B4EB5B5564A6ED7EA4D42856EFB4 - 1:0] IC2A6ECC367E2C82B97E73A57A8A79E1A ;
wire [I05264B2FA834FBEA729752C27B778963 - 1:0] I366D7D477BCE878309C2A4C6F4920631 ; wire I60B15FF62AA99717C8B7DA7D6912D281 ;
wire IA6BBDC90BCC6EF2E35BFA8D709343BF3 ; wire [I36A1B4EB5B5564A6ED7EA4D42856EFB4 - 1:0] I5631F39935597168A2C9D3656C66CB5C ;
wire [I6BAD12625217B36EDD0324B5AD4BB875 - 1:0] I1E2790529716BDA31237F724D6F3C1DA ; wire I8A3A10780386E36D927EC523D63F0852 ;
wire I366EB0B781FD462E1BDC374519E76C20 ; wire [I05F95435FA8D508B4820D9E064382614 - 1:0] I2CA1A324143051A0AFDEFB54659C657C ;
wire I704831C7406B6F1F8F643A5A69CA283F ; wire IA9BFFFC53E33C8CC8A916546D023AA92 ; wire [9:0] I68F165DF932475EADE453095B18725C5 ;
wire I4AE98FF3DA4D5A5EE68F8A14D9D781F4 ; wire IA5B2934FB33191AB00E5C1593870B4B4 ; wire [I64BB723AC8F87F7AEBA73BF190ED5F8F
- 1:0] I847247D81806836A31E3F617617623A1 ;  assign ID7FCE45A65ADDB17F91F73A1B506BB5B = I366D7D477BCE878309C2A4C6F4920631 ;
assign I125028C7446331521D0434C10E8B0007 = I847247D81806836A31E3F617617623A1 ; assign I8BB939FF2AFDE7B2A1E480DCB61CE354
= I60B15FF62AA99717C8B7DA7D6912D281 ; assign IC9DE8233C6B1ADF4418EEF5B1F14BE49 = IA5B2934FB33191AB00E5C1593870B4B4 ;
assign I585F74DE05DD9C1C7070D6B4F6E181C2 = IA6BBDC90BCC6EF2E35BFA8D709343BF3 ; assign I233E0C0C8E5150F0CD8258F276D93942
= I1E2790529716BDA31237F724D6F3C1DA ; assign IBE0D6810EBD63B5C428623C578CF6D3A = I366EB0B781FD462E1BDC374519E76C20 ;
 assign {IA5B2934FB33191AB00E5C1593870B4B4 , I847247D81806836A31E3F617617623A1 } = I2CA1A324143051A0AFDEFB54659C657C ;
assign I4AE98FF3DA4D5A5EE68F8A14D9D781F4 = ~I9ED2A9117D3AEAF54CBA7AD69083BCB7 ; generate if (IFA55551D85BC21F7BB69A4B7EF5E7D87
== 1) begin assign I704831C7406B6F1F8F643A5A69CA283F = I2CA1A324143051A0AFDEFB54659C657C [29]; assign IA9BFFFC53E33C8CC8A916546D023AA92
= I2CA1A324143051A0AFDEFB54659C657C [30]; assign I68F165DF932475EADE453095B18725C5 = I2CA1A324143051A0AFDEFB54659C657C [9:0];
end else begin assign I704831C7406B6F1F8F643A5A69CA283F = I2CA1A324143051A0AFDEFB54659C657C [61]; assign IA9BFFFC53E33C8CC8A916546D023AA92
= I2CA1A324143051A0AFDEFB54659C657C [62]; assign I68F165DF932475EADE453095B18725C5 = I2CA1A324143051A0AFDEFB54659C657C [41:32];
end endgenerate  IA8C351750B9DBEE4D8ADA94748C8E5D1 #( .I61D0345D311EC6FFC08DDDECE5F6127A (IB71844FFA3AB85FEF45EAB4D35395752 ),
.I5C6C6CD7723900C21B3A76E887CEE164 (I5C6C6CD7723900C21B3A76E887CEE164 ), .I64BB723AC8F87F7AEBA73BF190ED5F8F (I64BB723AC8F87F7AEBA73BF190ED5F8F )
) IB420C4D1279F971E867FA537CA4D6E82 ( .I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .ICCFB0F435B37370076102F325BC08D20
(ICCFB0F435B37370076102F325BC08D20 ), .I8F36BEAA79ADAC31FBCBAC1B805C772E (I704831C7406B6F1F8F643A5A69CA283F ), .IE52544EAEF6757A8A982FC14CE507F8C
(IA9BFFFC53E33C8CC8A916546D023AA92 ), .IAC8BFFA8C250FC35278EA36BA7C00B42 (I68F165DF932475EADE453095B18725C5 ), .I27CF4DD7FCBC7E0A229344EDF94F2651
(I27CF4DD7FCBC7E0A229344EDF94F2651 ), .I1A55EB74BDB9184AA980B07905C85479 (I1A55EB74BDB9184AA980B07905C85479 ), .IC79EC9A9F373F4B71374BDF6EDD31DE6
(1'b0), .ID8853B025150C80EE45BBA98E5BEA3A8 (I48D61F5A0B5732A58912433B42CD9D0C ), .I04BC24D2B6403E54A64DE9E6C9ABAA2B
(I04BC24D2B6403E54A64DE9E6C9ABAA2B ), .I3F6FB755DC9826D564C143FF9E32F032 (I3F6FB755DC9826D564C143FF9E32F032 ), .IE315CDCA06C9620D5C0AB966E553F0C3
(IE315CDCA06C9620D5C0AB966E553F0C3 ), .I7740E93179670969593F64CBA98864D9 (IC2A6ECC367E2C82B97E73A57A8A79E1A ), .I89011D8BA1FC92A73CD875E098FE685C
(I5631F39935597168A2C9D3656C66CB5C ), .I7D649F765882BD862315E777ABA5263F (IFAF7F03355554E59A3861F8A72D71CA5 ), .I87AD4A36141619A102AD5166323D80AB
(I8A3A10780386E36D927EC523D63F0852 ), .ID7FCE45A65ADDB17F91F73A1B506BB5B (I366D7D477BCE878309C2A4C6F4920631 ), .I8BB939FF2AFDE7B2A1E480DCB61CE354
(I60B15FF62AA99717C8B7DA7D6912D281 ), .I585F74DE05DD9C1C7070D6B4F6E181C2 (IA6BBDC90BCC6EF2E35BFA8D709343BF3 ), .I233E0C0C8E5150F0CD8258F276D93942
(I1E2790529716BDA31237F724D6F3C1DA ), .IBE0D6810EBD63B5C428623C578CF6D3A (I366EB0B781FD462E1BDC374519E76C20 ) );
pmi_ram_dp # ( .pmi_wr_addr_depth (IB71844FFA3AB85FEF45EAB4D35395752 ), .pmi_wr_addr_width (I36A1B4EB5B5564A6ED7EA4D42856EFB4 ),
.pmi_wr_data_width (I05F95435FA8D508B4820D9E064382614 ), .pmi_rd_addr_depth (IB71844FFA3AB85FEF45EAB4D35395752 ),
.pmi_rd_addr_width (I36A1B4EB5B5564A6ED7EA4D42856EFB4 ), .pmi_rd_data_width (I05F95435FA8D508B4820D9E064382614 ),
.pmi_regmode ("reg"), .pmi_family (I66C185998F46A7148163982E39BCD296 ), .module_type ("pmi_ram_dp") ) I32900CECD80193336B4F376406D5DFF6
( .Data (IFAF7F03355554E59A3861F8A72D71CA5 ), .RdAddress (IC2A6ECC367E2C82B97E73A57A8A79E1A ), .RdClockEn (1'b1),
.RdClock (ICCFB0F435B37370076102F325BC08D20 ), .Reset (I4AE98FF3DA4D5A5EE68F8A14D9D781F4 ), .WE (I8A3A10780386E36D927EC523D63F0852 ),
.WrAddress (I5631F39935597168A2C9D3656C66CB5C ), .WrClockEn (1'b1), .WrClock (ICCFB0F435B37370076102F325BC08D20 ),
.Q (I2CA1A324143051A0AFDEFB54659C657C ) ); endmodule 
  module I8489B3291801D4F3BE8AED05E26C4566 #( parameter I87C69AEB153025D890F0A7CE399F00FE = 2 ) ( input wire ICCFB0F435B37370076102F325BC08D20 ,
input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire [12:0] I488999E90FEFB5E25518723EB6105532 , input wire
[8:0] IB064E00468F70C38840D1D271524C6C8 , input wire [12:0] IE4E19EA6F3F828B3B44ED1E4D36558F7 , input wire [8:0]
I537C738B170D60A42A1F6FDA4547BACC , input wire [12:0] IA29842BA67669CD8D75483E633C363F0 , input wire [8:0] IB9E3BDBEE7C442BA69CD12711DA40F71 ,
input wire IABD5FBD9A9966396ACABECC997D287C6 , input wire I06326CB6C7B31C2BC01AEF85D6548C61 , input wire IADC13C79970748AA5DA1B07EC1C4290D ,
input wire ICDFC5D4FA0C2CE90CDF9381D077D8CE2 , input wire I756CF2AA8135461091FB5662DDE3111E , input wire [31:0]
I2687BB96A4E1D15035B283D3FDF616CC , input wire [31:0] I2EF8304B3AEA32E6C6F568223FAD9CBA , input wire [31:0] I369C6CA451B73B45E1F8D4D8AA53C2AD ,
input wire [31:0] IE81278F89BAA90C1F6EF0784D0DE2F62 , input wire I2F86B5F8620848A51ED4F1F736CF8825 , input wire
I63FDDFAA5AB093F3BB343A8C133F3BAF , input wire IE7F8A35B24BC8805CAD86FD378C18296 , input wire IAB90D3559ED5004EBCCD9D73A2928E3F ,
input wire [I87C69AEB153025D890F0A7CE399F00FE - 1:0] I75EB9BE30F2D20C56659251E3B505209 , input wire I3E8F0524CDEE96F573376A6BF670184B ,
input wire I17066520A25539E7F98555DFF7832BBE , output wire [15:0] IB33B8D629A269D1BC3D79902EE2EB312 , output wire
I4A4976CAF016EA789DCDB7AA131246C3 , output wire I5ADFC7E7F8B570F5258C2813D0020950 , output wire I1FD27F5D298FA5493F3F510610F19E4E ,
output wire ID7F4713F32DABD57E54222A946FA802F , output wire IADE62F3832E7DA9091E0F5B2EBC50F9C , output wire I3443654006276E8DC7EE67AAE2283C64 ,
output wire I4FD27244D7DB92B0548A7AE35BDEDE28 , output wire IDB44E9A441DC017FFA044AB8E232791F ); `include "tlp_qcodes.v"
localparam IC8B5868CE6CCCFF479B9D42AE258A6C9 = 4'b0000, IE52A4905856745CF06589D8BBCBF62C0 = 4'b0001, I797FF78A781B011D1491E42DA6E8E636
= 4'b0010, I1829FA88EF5AD31D47831CE2250D10F7 = 4'b0011, I2F1344D3FD89FDF0D046D2CFE8B81756 = 4'b0100, I81433A6080C7D6A889CE2862E42D5F2C
= 4'b0101, IFCC4638207CC2B4943B7A3D236493B68 = 4'b0110, I60218F936AC6C7F041F5C51CF271A588 = 4'b0111, I819A59AEE1BB0A106C574B93C030EA0A
= 4'b1000, I4B14F35045D0C6D4ACC52F05548C8ED0 = 4'b1001, I805E1EB4F502A27328E7ED208D7524F0 = 4'b1010, IB63534807AE73A9DD6F73F942EAAB356
= 4'b1011;  reg [12:0] I31C96A05CDA83684954EE47D715D4665 ; reg [12:0] I8E17DAB6BBC782E384ABBDDC296D791C ; reg I3565B787C28964F625269B34EE86A5CA ;
reg IDA82F4C78A43B62E1C09ED19A1443221 ; reg IF4B2F356412545C21578876129150C2F ; reg [1:0] I094BDF55C12CD5E2524B36CC933CFAE3 ;
reg I36AB316E2312154193B60465E4A46981 ; reg [1:0] IF3BFEFDD423F2FF0D209290C782C2472 ; reg [10:0] IF8163AD5BD15021B831D22F3FD61BA6A ;
reg [15:0] IE5C1CB646B621DD5D037AA5F5961D901 ; reg I23A5651CB59E99C9EF06BE735CE54321 ; reg I9B1524315BD1F28EE8423E6A4D5CA375 ;
reg I042EEC1DF7AD7810D40B515154D92853 ; reg [31:0] ID0A5ECECBEC8CE692F380DDF069E842F ; reg [31:0] IBC3E292376641E5290114F38B65B8702 ;
reg ICE47914C96690A70DF3F7A7C01052696 ; reg I0AAA85DA619AFA12BBAB9F4AF77B9C6C ; reg IB27F7D37271B47673F001712E52E16F2 ;
reg IDD78F0F33DD4EEA1A7F1111B4B04E3EF ; reg I41D6A7D674F63A59E5DBBE00AA282E14 ; reg I23B9845BB3A093CE647D68158F400F36 ;
reg I9542E55FC3D72D91960B79EC50367A55 ; reg I0CA51557A90D8B4060C406DC652C2485 ; reg [10:0] I28BEA4229042F20DC4BAC5A80E0CF354 ;
reg I57700DAA2CEC60C16029DE31DBC7F36B ; reg I6513C757AD9B98D491547EBB8D69BC7D ; reg I297D3FE7B056FB743893BCFC1B67D805 ;
reg I4F5985BF6243B7F0468BA4DD2B5D2E06 ; reg [IC7701945BBBE654661A8C2F153881F63 :0] I91A6742D4BEEA347CB6EDF3386EC70F6 ;
reg IE3F232999F09A0949531BDA44AC0700A ; reg [3:0] I569BD691A4BB295D836212F3738D46B4 ; reg [3:0] IFC499732997C1DCC89CB1F5E9F9C4CB3 ;
wire I62AEDB14F0B7669ACCEF627D809BAF73 ; wire I7EAA8AFFB2BC9D190B3626833AF5EBD8 ;  assign IB33B8D629A269D1BC3D79902EE2EB312
= IE5C1CB646B621DD5D037AA5F5961D901 ; assign I4A4976CAF016EA789DCDB7AA131246C3 = I23A5651CB59E99C9EF06BE735CE54321 ;
assign I5ADFC7E7F8B570F5258C2813D0020950 = (I569BD691A4BB295D836212F3738D46B4 == I60218F936AC6C7F041F5C51CF271A588 )
? 1'b1 : 1'b0; assign I1FD27F5D298FA5493F3F510610F19E4E = I9B1524315BD1F28EE8423E6A4D5CA375 ; assign ID7F4713F32DABD57E54222A946FA802F
= ICE47914C96690A70DF3F7A7C01052696 ; assign IADE62F3832E7DA9091E0F5B2EBC50F9C = I0AAA85DA619AFA12BBAB9F4AF77B9C6C ;
assign I3443654006276E8DC7EE67AAE2283C64 = IB27F7D37271B47673F001712E52E16F2 ; assign I4FD27244D7DB92B0548A7AE35BDEDE28
= IDD78F0F33DD4EEA1A7F1111B4B04E3EF ; assign IDB44E9A441DC017FFA044AB8E232791F = (I569BD691A4BB295D836212F3738D46B4
== IE52A4905856745CF06589D8BBCBF62C0 ) ? 1'b1 : 1'b0;  assign I62AEDB14F0B7669ACCEF627D809BAF73 = ICE47914C96690A70DF3F7A7C01052696
| I0AAA85DA619AFA12BBAB9F4AF77B9C6C | IB27F7D37271B47673F001712E52E16F2 | IDD78F0F33DD4EEA1A7F1111B4B04E3EF ; assign
I7EAA8AFFB2BC9D190B3626833AF5EBD8 = I06326CB6C7B31C2BC01AEF85D6548C61 | IADC13C79970748AA5DA1B07EC1C4290D | ICDFC5D4FA0C2CE90CDF9381D077D8CE2
| I756CF2AA8135461091FB5662DDE3111E ;  always @(*) begin IFC499732997C1DCC89CB1F5E9F9C4CB3 = I569BD691A4BB295D836212F3738D46B4 ;
case (I569BD691A4BB295D836212F3738D46B4 ) IC8B5868CE6CCCFF479B9D42AE258A6C9 : begin if (~I3E8F0524CDEE96F573376A6BF670184B )
IFC499732997C1DCC89CB1F5E9F9C4CB3 = IE52A4905856745CF06589D8BBCBF62C0 ; end IE52A4905856745CF06589D8BBCBF62C0 :
begin IFC499732997C1DCC89CB1F5E9F9C4CB3 = I797FF78A781B011D1491E42DA6E8E636 ; end I797FF78A781B011D1491E42DA6E8E636
: begin if (I17066520A25539E7F98555DFF7832BBE == 1'b1) IFC499732997C1DCC89CB1F5E9F9C4CB3 = I1829FA88EF5AD31D47831CE2250D10F7 ;
end I1829FA88EF5AD31D47831CE2250D10F7 : begin IFC499732997C1DCC89CB1F5E9F9C4CB3 = I2F1344D3FD89FDF0D046D2CFE8B81756 ;
end I2F1344D3FD89FDF0D046D2CFE8B81756 : begin IFC499732997C1DCC89CB1F5E9F9C4CB3 = I81433A6080C7D6A889CE2862E42D5F2C ;
end I81433A6080C7D6A889CE2862E42D5F2C : begin if (I7EAA8AFFB2BC9D190B3626833AF5EBD8 ) IFC499732997C1DCC89CB1F5E9F9C4CB3
= IFCC4638207CC2B4943B7A3D236493B68 ; end IFCC4638207CC2B4943B7A3D236493B68 : begin if (I3565B787C28964F625269B34EE86A5CA )
IFC499732997C1DCC89CB1F5E9F9C4CB3 = I60218F936AC6C7F041F5C51CF271A588 ; end I60218F936AC6C7F041F5C51CF271A588 :
begin if (IABD5FBD9A9966396ACABECC997D287C6 ) IFC499732997C1DCC89CB1F5E9F9C4CB3 = I819A59AEE1BB0A106C574B93C030EA0A ;
end I819A59AEE1BB0A106C574B93C030EA0A : begin IFC499732997C1DCC89CB1F5E9F9C4CB3 = I4B14F35045D0C6D4ACC52F05548C8ED0 ;
end I4B14F35045D0C6D4ACC52F05548C8ED0 : begin IFC499732997C1DCC89CB1F5E9F9C4CB3 = I805E1EB4F502A27328E7ED208D7524F0 ;
end I805E1EB4F502A27328E7ED208D7524F0 : begin if (IE3F232999F09A0949531BDA44AC0700A == 1'b1) if (I23A5651CB59E99C9EF06BE735CE54321
== 1'b1) IFC499732997C1DCC89CB1F5E9F9C4CB3 = IC8B5868CE6CCCFF479B9D42AE258A6C9 ; else begin if (IF3BFEFDD423F2FF0D209290C782C2472
== 0) IFC499732997C1DCC89CB1F5E9F9C4CB3 = IB63534807AE73A9DD6F73F942EAAB356 ; end end IB63534807AE73A9DD6F73F942EAAB356
: begin if (I23A5651CB59E99C9EF06BE735CE54321 == 1'b1) IFC499732997C1DCC89CB1F5E9F9C4CB3 = IC8B5868CE6CCCFF479B9D42AE258A6C9 ;
end default : begin end endcase end  always @(*) begin case (I91A6742D4BEEA347CB6EDF3386EC70F6 ) I83EA49D19551ED8C672BF332D148F920
: begin IBC3E292376641E5290114F38B65B8702 = I2687BB96A4E1D15035B283D3FDF616CC ; end I373604D502FD927695BB13BAA1D3443F
: begin IBC3E292376641E5290114F38B65B8702 = I2EF8304B3AEA32E6C6F568223FAD9CBA ; end IA687834EBB97378F700DB12C9394F09F
: begin IBC3E292376641E5290114F38B65B8702 = I369C6CA451B73B45E1F8D4D8AA53C2AD ; end IF59ACE7A9B4E430EAAD83B6808CA927D
: begin IBC3E292376641E5290114F38B65B8702 = IE81278F89BAA90C1F6EF0784D0DE2F62 ; end endcase end  always @(posedge
ICCFB0F435B37370076102F325BC08D20 or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin if (~I9ED2A9117D3AEAF54CBA7AD69083BCB7 )
begin I31C96A05CDA83684954EE47D715D4665 <= 13'b0; I8E17DAB6BBC782E384ABBDDC296D791C <= 13'b0; I3565B787C28964F625269B34EE86A5CA
<= 1'b0; IDA82F4C78A43B62E1C09ED19A1443221 <= 1'b0; IF4B2F356412545C21578876129150C2F <= 1'b0; I094BDF55C12CD5E2524B36CC933CFAE3
<= 2'b0; I36AB316E2312154193B60465E4A46981 <= 1'b1; IF3BFEFDD423F2FF0D209290C782C2472 <= 10'b0; IF8163AD5BD15021B831D22F3FD61BA6A
<= 10'b0; IE5C1CB646B621DD5D037AA5F5961D901 <= 16'b0; I23A5651CB59E99C9EF06BE735CE54321 <= 1'b0; I9B1524315BD1F28EE8423E6A4D5CA375
<= 1'b0; I042EEC1DF7AD7810D40B515154D92853 <= 1'b0; ICE47914C96690A70DF3F7A7C01052696 <= 1'b0; I0AAA85DA619AFA12BBAB9F4AF77B9C6C
<= 1'b0; IB27F7D37271B47673F001712E52E16F2 <= 1'b0; IDD78F0F33DD4EEA1A7F1111B4B04E3EF <= 1'b0; I41D6A7D674F63A59E5DBBE00AA282E14
<= 1'b0; I23B9845BB3A093CE647D68158F400F36 <= 1'b0; I9542E55FC3D72D91960B79EC50367A55 <= 1'b0; I0CA51557A90D8B4060C406DC652C2485
<= 1'b0; I28BEA4229042F20DC4BAC5A80E0CF354 <= 10'b0; I57700DAA2CEC60C16029DE31DBC7F36B <= 1'b1; I6513C757AD9B98D491547EBB8D69BC7D
<= 1'b0; I297D3FE7B056FB743893BCFC1B67D805 <= 1'b0; I4F5985BF6243B7F0468BA4DD2B5D2E06 <= 1'b0; I91A6742D4BEEA347CB6EDF3386EC70F6
<= 2'b0; I569BD691A4BB295D836212F3738D46B4 <= IC8B5868CE6CCCFF479B9D42AE258A6C9 ; IE3F232999F09A0949531BDA44AC0700A
<= 1'b0; end else begin I31C96A05CDA83684954EE47D715D4665 <= I488999E90FEFB5E25518723EB6105532 ; I8E17DAB6BBC782E384ABBDDC296D791C
<= IA29842BA67669CD8D75483E633C363F0 ; I23A5651CB59E99C9EF06BE735CE54321 <= 1'b0; I9B1524315BD1F28EE8423E6A4D5CA375
<= 1'b0; I042EEC1DF7AD7810D40B515154D92853 <= ICE47914C96690A70DF3F7A7C01052696 | I0AAA85DA619AFA12BBAB9F4AF77B9C6C
| IB27F7D37271B47673F001712E52E16F2 | IDD78F0F33DD4EEA1A7F1111B4B04E3EF ; ICE47914C96690A70DF3F7A7C01052696 <= 1'b0;
I0AAA85DA619AFA12BBAB9F4AF77B9C6C <= 1'b0; IB27F7D37271B47673F001712E52E16F2 <= 1'b0; IDD78F0F33DD4EEA1A7F1111B4B04E3EF
<= 1'b0; I41D6A7D674F63A59E5DBBE00AA282E14 <= ~I2F86B5F8620848A51ED4F1F736CF8825 ; I23B9845BB3A093CE647D68158F400F36
<= ~I63FDDFAA5AB093F3BB343A8C133F3BAF ; I9542E55FC3D72D91960B79EC50367A55 <= ~IE7F8A35B24BC8805CAD86FD378C18296 ;
I0CA51557A90D8B4060C406DC652C2485 <= ~IAB90D3559ED5004EBCCD9D73A2928E3F ; I6513C757AD9B98D491547EBB8D69BC7D <= (ID0A5ECECBEC8CE692F380DDF069E842F [1:0]
== 2'b0) ? ((I31C96A05CDA83684954EE47D715D4665 >= ID0A5ECECBEC8CE692F380DDF069E842F [9:2]) ? I41D6A7D674F63A59E5DBBE00AA282E14
: 1'b0) : ((I31C96A05CDA83684954EE47D715D4665 > ID0A5ECECBEC8CE692F380DDF069E842F [9:2]) ? I41D6A7D674F63A59E5DBBE00AA282E14
: 1'b0); I297D3FE7B056FB743893BCFC1B67D805 <= (ID0A5ECECBEC8CE692F380DDF069E842F [1:0] == 2'b0) ? ((I8E17DAB6BBC782E384ABBDDC296D791C
>= ID0A5ECECBEC8CE692F380DDF069E842F [9:2]) ? I9542E55FC3D72D91960B79EC50367A55 : 1'b0) : ((I8E17DAB6BBC782E384ABBDDC296D791C
> ID0A5ECECBEC8CE692F380DDF069E842F [9:2]) ? I9542E55FC3D72D91960B79EC50367A55 : 1'b0); I4F5985BF6243B7F0468BA4DD2B5D2E06
<= (ID0A5ECECBEC8CE692F380DDF069E842F [1:0] == 2'b0) ? ((I8E17DAB6BBC782E384ABBDDC296D791C >= ID0A5ECECBEC8CE692F380DDF069E842F [9:2])
? I0CA51557A90D8B4060C406DC652C2485 : 1'b0) : ((I8E17DAB6BBC782E384ABBDDC296D791C > ID0A5ECECBEC8CE692F380DDF069E842F [9:2])
? I0CA51557A90D8B4060C406DC652C2485 : 1'b0); I569BD691A4BB295D836212F3738D46B4 <= IFC499732997C1DCC89CB1F5E9F9C4CB3 ;
IE3F232999F09A0949531BDA44AC0700A <= I7EAA8AFFB2BC9D190B3626833AF5EBD8 ; if (I62AEDB14F0B7669ACCEF627D809BAF73 ==
1'b1) begin if (I094BDF55C12CD5E2524B36CC933CFAE3 > 0) begin I094BDF55C12CD5E2524B36CC933CFAE3 <= I094BDF55C12CD5E2524B36CC933CFAE3
- 1; I36AB316E2312154193B60465E4A46981 <= (I094BDF55C12CD5E2524B36CC933CFAE3 == 1) ? 1'b1 : 1'b0; end else if (I28BEA4229042F20DC4BAC5A80E0CF354
> 0) begin I28BEA4229042F20DC4BAC5A80E0CF354 <= I28BEA4229042F20DC4BAC5A80E0CF354 - 1; I57700DAA2CEC60C16029DE31DBC7F36B
<= (I28BEA4229042F20DC4BAC5A80E0CF354 == 1) ? 1'b1 : 1'b0; end end if (I17066520A25539E7F98555DFF7832BBE == 1'b1)
I91A6742D4BEEA347CB6EDF3386EC70F6 <= I75EB9BE30F2D20C56659251E3B505209 ; if (I042EEC1DF7AD7810D40B515154D92853 ==
1'b1) case (I91A6742D4BEEA347CB6EDF3386EC70F6 ) I83EA49D19551ED8C672BF332D148F920 : ID0A5ECECBEC8CE692F380DDF069E842F
<= I2687BB96A4E1D15035B283D3FDF616CC ; I373604D502FD927695BB13BAA1D3443F : ID0A5ECECBEC8CE692F380DDF069E842F <=
I2EF8304B3AEA32E6C6F568223FAD9CBA ; IA687834EBB97378F700DB12C9394F09F : ID0A5ECECBEC8CE692F380DDF069E842F <= I369C6CA451B73B45E1F8D4D8AA53C2AD ;
IF59ACE7A9B4E430EAAD83B6808CA927D : ID0A5ECECBEC8CE692F380DDF069E842F <= IE81278F89BAA90C1F6EF0784D0DE2F62 ; default
: begin end endcase case (I569BD691A4BB295D836212F3738D46B4 ) IE52A4905856745CF06589D8BBCBF62C0 : begin I3565B787C28964F625269B34EE86A5CA
<= 1'b0; end I1829FA88EF5AD31D47831CE2250D10F7 : begin ICE47914C96690A70DF3F7A7C01052696 <= (I91A6742D4BEEA347CB6EDF3386EC70F6
== I83EA49D19551ED8C672BF332D148F920 ) ? 1'b1 : 1'b0; I0AAA85DA619AFA12BBAB9F4AF77B9C6C <= (I91A6742D4BEEA347CB6EDF3386EC70F6
== I373604D502FD927695BB13BAA1D3443F ) ? 1'b1 : 1'b0; IB27F7D37271B47673F001712E52E16F2 <= (I91A6742D4BEEA347CB6EDF3386EC70F6
== IA687834EBB97378F700DB12C9394F09F ) ? 1'b1 : 1'b0; IDD78F0F33DD4EEA1A7F1111B4B04E3EF <= (I91A6742D4BEEA347CB6EDF3386EC70F6
== IF59ACE7A9B4E430EAAD83B6808CA927D ) ? 1'b1 : 1'b0; end I2F1344D3FD89FDF0D046D2CFE8B81756 : begin end I81433A6080C7D6A889CE2862E42D5F2C
: begin if (I042EEC1DF7AD7810D40B515154D92853 == 1'b0) begin IDA82F4C78A43B62E1C09ED19A1443221 <= ((I91A6742D4BEEA347CB6EDF3386EC70F6
== I83EA49D19551ED8C672BF332D148F920 ) || (I91A6742D4BEEA347CB6EDF3386EC70F6 == IA687834EBB97378F700DB12C9394F09F )
|| (I91A6742D4BEEA347CB6EDF3386EC70F6 == IF59ACE7A9B4E430EAAD83B6808CA927D )) ? ID0A5ECECBEC8CE692F380DDF069E842F [30]
: 1'b0; IF4B2F356412545C21578876129150C2F <= ((I91A6742D4BEEA347CB6EDF3386EC70F6 == I373604D502FD927695BB13BAA1D3443F )
|| (I91A6742D4BEEA347CB6EDF3386EC70F6 == IA687834EBB97378F700DB12C9394F09F ) || (I91A6742D4BEEA347CB6EDF3386EC70F6
== IF59ACE7A9B4E430EAAD83B6808CA927D )) ? ID0A5ECECBEC8CE692F380DDF069E842F [29] : 1'b0; end end IFCC4638207CC2B4943B7A3D236493B68
: begin I36AB316E2312154193B60465E4A46981 <= 1'b0; IF8163AD5BD15021B831D22F3FD61BA6A <= ID0A5ECECBEC8CE692F380DDF069E842F [9:0];
I28BEA4229042F20DC4BAC5A80E0CF354 <= (IDA82F4C78A43B62E1C09ED19A1443221 == 1'b1) ? ID0A5ECECBEC8CE692F380DDF069E842F [9:0]
: 10'b0; I57700DAA2CEC60C16029DE31DBC7F36B <= ~IDA82F4C78A43B62E1C09ED19A1443221 ;  if (IF4B2F356412545C21578876129150C2F )
begin I094BDF55C12CD5E2524B36CC933CFAE3 <= 2'b11; IF3BFEFDD423F2FF0D209290C782C2472 <= 2'b10; end else begin I094BDF55C12CD5E2524B36CC933CFAE3
<= 2'b10; IF3BFEFDD423F2FF0D209290C782C2472 <= 2'b01; end case (I91A6742D4BEEA347CB6EDF3386EC70F6 ) I83EA49D19551ED8C672BF332D148F920
: begin if (IDA82F4C78A43B62E1C09ED19A1443221 ) I3565B787C28964F625269B34EE86A5CA <= (|IB064E00468F70C38840D1D271524C6C8 )
? I6513C757AD9B98D491547EBB8D69BC7D : 1'b0; else I3565B787C28964F625269B34EE86A5CA <= (|IB064E00468F70C38840D1D271524C6C8 )
? 1'b1 : 1'b0; end I373604D502FD927695BB13BAA1D3443F : begin I3565B787C28964F625269B34EE86A5CA <= (|I537C738B170D60A42A1F6FDA4547BACC )
? 1'b1 : 1'b0; end IA687834EBB97378F700DB12C9394F09F : begin if (IDA82F4C78A43B62E1C09ED19A1443221 ) I3565B787C28964F625269B34EE86A5CA
<= (|IB9E3BDBEE7C442BA69CD12711DA40F71 ) ? I297D3FE7B056FB743893BCFC1B67D805 : 1'b0; else I3565B787C28964F625269B34EE86A5CA
<= (|IB9E3BDBEE7C442BA69CD12711DA40F71 ) ? 1'b1 : 1'b0; end IF59ACE7A9B4E430EAAD83B6808CA927D : begin if (IDA82F4C78A43B62E1C09ED19A1443221 )
I3565B787C28964F625269B34EE86A5CA <= (|IB9E3BDBEE7C442BA69CD12711DA40F71 ) ? I4F5985BF6243B7F0468BA4DD2B5D2E06 :
1'b0; else I3565B787C28964F625269B34EE86A5CA <= (|IB9E3BDBEE7C442BA69CD12711DA40F71 ) ? 1'b1 : 1'b0; end endcase
end I60218F936AC6C7F041F5C51CF271A588 : begin IE5C1CB646B621DD5D037AA5F5961D901 <= (IABD5FBD9A9966396ACABECC997D287C6
== 1'b1) ? ID0A5ECECBEC8CE692F380DDF069E842F [31:16] : 16'b0; I9B1524315BD1F28EE8423E6A4D5CA375 <= IABD5FBD9A9966396ACABECC997D287C6 ;
ICE47914C96690A70DF3F7A7C01052696 <= (I91A6742D4BEEA347CB6EDF3386EC70F6 == I83EA49D19551ED8C672BF332D148F920 ) ?
IABD5FBD9A9966396ACABECC997D287C6 : 1'b0; I0AAA85DA619AFA12BBAB9F4AF77B9C6C <= (I91A6742D4BEEA347CB6EDF3386EC70F6
== I373604D502FD927695BB13BAA1D3443F ) ? IABD5FBD9A9966396ACABECC997D287C6 : 1'b0; IB27F7D37271B47673F001712E52E16F2
<= (I91A6742D4BEEA347CB6EDF3386EC70F6 == IA687834EBB97378F700DB12C9394F09F ) ? IABD5FBD9A9966396ACABECC997D287C6
: 1'b0; IDD78F0F33DD4EEA1A7F1111B4B04E3EF <= (I91A6742D4BEEA347CB6EDF3386EC70F6 == IF59ACE7A9B4E430EAAD83B6808CA927D )
? IABD5FBD9A9966396ACABECC997D287C6 : 1'b0; end I819A59AEE1BB0A106C574B93C030EA0A : begin IE5C1CB646B621DD5D037AA5F5961D901
<= (IABD5FBD9A9966396ACABECC997D287C6 == 1'b1) ? ID0A5ECECBEC8CE692F380DDF069E842F [15:0] : 16'b0; end I4B14F35045D0C6D4ACC52F05548C8ED0
: begin IE5C1CB646B621DD5D037AA5F5961D901 <= IBC3E292376641E5290114F38B65B8702 [31:16]; ICE47914C96690A70DF3F7A7C01052696
<= (I91A6742D4BEEA347CB6EDF3386EC70F6 == I83EA49D19551ED8C672BF332D148F920 ) ? 1'b1 : 1'b0; I0AAA85DA619AFA12BBAB9F4AF77B9C6C
<= (I91A6742D4BEEA347CB6EDF3386EC70F6 == I373604D502FD927695BB13BAA1D3443F ) ? 1'b1 : 1'b0; IB27F7D37271B47673F001712E52E16F2
<= (I91A6742D4BEEA347CB6EDF3386EC70F6 == IA687834EBB97378F700DB12C9394F09F ) ? 1'b1 : 1'b0; IDD78F0F33DD4EEA1A7F1111B4B04E3EF
<= (I91A6742D4BEEA347CB6EDF3386EC70F6 == IF59ACE7A9B4E430EAAD83B6808CA927D ) ? 1'b1 : 1'b0; end I805E1EB4F502A27328E7ED208D7524F0
: begin ICE47914C96690A70DF3F7A7C01052696 <= (I91A6742D4BEEA347CB6EDF3386EC70F6 == I83EA49D19551ED8C672BF332D148F920 )
? ~ICE47914C96690A70DF3F7A7C01052696 & (~I36AB316E2312154193B60465E4A46981 | (IDA82F4C78A43B62E1C09ED19A1443221
& ~I57700DAA2CEC60C16029DE31DBC7F36B )) : 1'b0; I0AAA85DA619AFA12BBAB9F4AF77B9C6C <= (I91A6742D4BEEA347CB6EDF3386EC70F6
== I373604D502FD927695BB13BAA1D3443F ) ? (~I0AAA85DA619AFA12BBAB9F4AF77B9C6C & ~I36AB316E2312154193B60465E4A46981 )
: 1'b0; IB27F7D37271B47673F001712E52E16F2 <= (I91A6742D4BEEA347CB6EDF3386EC70F6 == IA687834EBB97378F700DB12C9394F09F )
? ~IB27F7D37271B47673F001712E52E16F2 & (~I36AB316E2312154193B60465E4A46981 | (IDA82F4C78A43B62E1C09ED19A1443221
& ~I57700DAA2CEC60C16029DE31DBC7F36B )) : 1'b0; IDD78F0F33DD4EEA1A7F1111B4B04E3EF <= (I91A6742D4BEEA347CB6EDF3386EC70F6
== IF59ACE7A9B4E430EAAD83B6808CA927D ) ? (~IDD78F0F33DD4EEA1A7F1111B4B04E3EF & ~I57700DAA2CEC60C16029DE31DBC7F36B )
: 1'b0; if (IE3F232999F09A0949531BDA44AC0700A ) begin IF3BFEFDD423F2FF0D209290C782C2472 <= IF3BFEFDD423F2FF0D209290C782C2472
- 1; IE5C1CB646B621DD5D037AA5F5961D901 <= IBC3E292376641E5290114F38B65B8702 [31:16]; end else begin IE5C1CB646B621DD5D037AA5F5961D901
<= IBC3E292376641E5290114F38B65B8702 [15:0]; I23A5651CB59E99C9EF06BE735CE54321 <= ((IF3BFEFDD423F2FF0D209290C782C2472
== 0) && (IDA82F4C78A43B62E1C09ED19A1443221 == 1'b0)) ? 1'b1 : 1'b0; end end IB63534807AE73A9DD6F73F942EAAB356 :
begin ICE47914C96690A70DF3F7A7C01052696 <= (I91A6742D4BEEA347CB6EDF3386EC70F6 == I83EA49D19551ED8C672BF332D148F920 )
? (~ICE47914C96690A70DF3F7A7C01052696 & ~I57700DAA2CEC60C16029DE31DBC7F36B ) : 1'b0; IB27F7D37271B47673F001712E52E16F2
<= (I91A6742D4BEEA347CB6EDF3386EC70F6 == IA687834EBB97378F700DB12C9394F09F ) ? (~IB27F7D37271B47673F001712E52E16F2
& ~I57700DAA2CEC60C16029DE31DBC7F36B ) : 1'b0; IDD78F0F33DD4EEA1A7F1111B4B04E3EF <= (I91A6742D4BEEA347CB6EDF3386EC70F6
== IF59ACE7A9B4E430EAAD83B6808CA927D ) ? (~IDD78F0F33DD4EEA1A7F1111B4B04E3EF & ~I57700DAA2CEC60C16029DE31DBC7F36B )
: 1'b0; if (IE3F232999F09A0949531BDA44AC0700A ) begin IF8163AD5BD15021B831D22F3FD61BA6A <= IF8163AD5BD15021B831D22F3FD61BA6A
- 1; IE5C1CB646B621DD5D037AA5F5961D901 <= IBC3E292376641E5290114F38B65B8702 [31:16]; end else begin IE5C1CB646B621DD5D037AA5F5961D901
<= IBC3E292376641E5290114F38B65B8702 [15:0]; I23A5651CB59E99C9EF06BE735CE54321 <= (IF8163AD5BD15021B831D22F3FD61BA6A
== 1) ? I7EAA8AFFB2BC9D190B3626833AF5EBD8 : 1'b0; end end endcase end end endmodule 
  module I5AA57FA362D8C2F14DF19B01C99AE372 #( parameter I87C69AEB153025D890F0A7CE399F00FE = 2 ) ( input wire ICCFB0F435B37370076102F325BC08D20 ,
input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire [12:0] I488999E90FEFB5E25518723EB6105532 , input wire
[8:0] IB064E00468F70C38840D1D271524C6C8 , input wire [12:0] IE4E19EA6F3F828B3B44ED1E4D36558F7 , input wire [8:0]
I537C738B170D60A42A1F6FDA4547BACC , input wire [12:0] IA29842BA67669CD8D75483E633C363F0 , input wire [8:0] IB9E3BDBEE7C442BA69CD12711DA40F71 ,
input wire IABD5FBD9A9966396ACABECC997D287C6 , input wire IFCFFF8448F5E6821B40C6CEE3548693A , input wire [2:0] I5CE5D2469FD5560C1773C754FC1E0C4A ,
input wire ID965E2D89D1047516134A3EED50CB8AE , input wire IC4019EF7E804F3D95AAA442EFE259D86 , input wire I8488C49C8D5977759183D4580A2BF116 ,
input wire I029FEAF1B2BC1E56CC9E23C77E352703 , input wire IE4A11C65C530DD3B14BE1A05F3324401 , input wire I06326CB6C7B31C2BC01AEF85D6548C61 ,
input wire IADC13C79970748AA5DA1B07EC1C4290D , input wire ICDFC5D4FA0C2CE90CDF9381D077D8CE2 , input wire I756CF2AA8135461091FB5662DDE3111E ,
input wire [63:0] I2687BB96A4E1D15035B283D3FDF616CC , input wire [63:0] I2EF8304B3AEA32E6C6F568223FAD9CBA , input
wire [63:0] I369C6CA451B73B45E1F8D4D8AA53C2AD , input wire [63:0] IE81278F89BAA90C1F6EF0784D0DE2F62 , input wire
I2F86B5F8620848A51ED4F1F736CF8825 , input wire I63FDDFAA5AB093F3BB343A8C133F3BAF , input wire IE7F8A35B24BC8805CAD86FD378C18296 ,
input wire IAB90D3559ED5004EBCCD9D73A2928E3F , input wire [I87C69AEB153025D890F0A7CE399F00FE - 1:0] I75EB9BE30F2D20C56659251E3B505209 ,
input wire I3E8F0524CDEE96F573376A6BF670184B , input wire I17066520A25539E7F98555DFF7832BBE , output wire [63:0]
IB33B8D629A269D1BC3D79902EE2EB312 , output wire I1E494BBA2ECB063404DBB73667CC7E8D , output wire I4A4976CAF016EA789DCDB7AA131246C3 ,
output wire I5ADFC7E7F8B570F5258C2813D0020950 , output wire I1FD27F5D298FA5493F3F510610F19E4E , output wire [1:0]
IEA9D116BFADD4042E3D3AD0C618B652A , output wire I418D7ADEC09B065FFE6565D649D285B6 , output wire IF2B42773D268BA706D29FCCFCB799AF9 ,
output wire I470C1C74A2768E559679EE12280C8506 , output wire I513461A4DA46CAA79BEC76A8DE8E2A98 , output wire ID7F4713F32DABD57E54222A946FA802F ,
output wire IADE62F3832E7DA9091E0F5B2EBC50F9C , output wire I3443654006276E8DC7EE67AAE2283C64 , output wire I4FD27244D7DB92B0548A7AE35BDEDE28 ,
output wire IDB44E9A441DC017FFA044AB8E232791F ); `include "tlp_qcodes.v"
localparam IC8B5868CE6CCCFF479B9D42AE258A6C9 = 4'b0000, IE52A4905856745CF06589D8BBCBF62C0 = 4'b0001, I797FF78A781B011D1491E42DA6E8E636
= 4'b0010, I1829FA88EF5AD31D47831CE2250D10F7 = 4'b0011, IFCC4638207CC2B4943B7A3D236493B68 = 4'b0100, I60218F936AC6C7F041F5C51CF271A588
= 4'b0101, IB784FFF6C985E87492B9D6F18C3910AE = 4'b0110, I293F67166A255C4EDC66C70F19551F8E = 4'b0111, I4ACB8367D46F2FB66718F5798E1F145F
= 4'b1000;  reg [12:0] I31C96A05CDA83684954EE47D715D4665 ; reg [12:0] I8E17DAB6BBC782E384ABBDDC296D791C ; reg I3565B787C28964F625269B34EE86A5CA ;
reg IDA82F4C78A43B62E1C09ED19A1443221 ; reg IF4B2F356412545C21578876129150C2F ; reg I928068FFB24833BA6A7A11BA59B8E040 ;
reg [63:0] IE5C1CB646B621DD5D037AA5F5961D901 ; reg I1742675C5CD0344DCC6E13EC6252ED0A ; reg I23A5651CB59E99C9EF06BE735CE54321 ;
reg IA1961DC2B849519BBCB37762269BB321 ; reg I9B1524315BD1F28EE8423E6A4D5CA375 ; reg I9A1E8CC9229E6A5D88D5CD96FBFE935D ;
reg [2:0] I637157BC0B4BC09421F86528FA1C6F22 ; reg I4DF8AE19A28761F0B98980365AEA794E ; reg [1:0] I3C78D9AB59D6164851A819C5BA6C7C04 ;
reg IE12E3E0C53D89CE85C02DAFD3FB81244 ; reg I8D8CDA8F60D3F8D5F51CD56B899536F8 ; reg IC373345D0993637162B568673C9F7143 ;
reg I5EBE440016CA0416EE3C2682065DDD85 ; reg [63:0] IBC3E292376641E5290114F38B65B8702 ; reg [63:0] IAA1E53CD0AE56DE019EFC1482B0134D6 ;
reg [63:0] I202B51CA022B3340D53544DEDC73872F ; reg [63:0] I37215D983C07F0C522E39A48B1F83101 ; reg [63:0] I1F1327610E72511D7678CF70DE3685C6 ;
reg I68014B0A38604EDB8B664C2C5CD25C03 ; reg I41D6A7D674F63A59E5DBBE00AA282E14 ; reg I23B9845BB3A093CE647D68158F400F36 ;
reg I9542E55FC3D72D91960B79EC50367A55 ; reg I0CA51557A90D8B4060C406DC652C2485 ; reg [10:0] I28BEA4229042F20DC4BAC5A80E0CF354 ;
reg I6513C757AD9B98D491547EBB8D69BC7D ; reg I297D3FE7B056FB743893BCFC1B67D805 ; reg I4F5985BF6243B7F0468BA4DD2B5D2E06 ;
reg [IC7701945BBBE654661A8C2F153881F63 :0] I91A6742D4BEEA347CB6EDF3386EC70F6 ; reg [3:0] I569BD691A4BB295D836212F3738D46B4 ;
reg [3:0] IFC499732997C1DCC89CB1F5E9F9C4CB3 ; reg [2:0] I45917910AA4CC0F07BA1A8EF74FE6FEF ; wire ID59D28ABECF4E3544E08856EFCBC426D ;
wire IE31D0AF3EFB3124913CD965CEE542B24 ; wire IA21F6AD8A9BCF2140ECB6EE68E7A9FC5 ; wire I7EAA8AFFB2BC9D190B3626833AF5EBD8 ;
 assign IB33B8D629A269D1BC3D79902EE2EB312 = IE5C1CB646B621DD5D037AA5F5961D901 ; assign I1E494BBA2ECB063404DBB73667CC7E8D
= I1742675C5CD0344DCC6E13EC6252ED0A ; assign I4A4976CAF016EA789DCDB7AA131246C3 = I23A5651CB59E99C9EF06BE735CE54321 ;
assign I5ADFC7E7F8B570F5258C2813D0020950 = IA1961DC2B849519BBCB37762269BB321 ; assign I1FD27F5D298FA5493F3F510610F19E4E
= I9B1524315BD1F28EE8423E6A4D5CA375 ; assign IEA9D116BFADD4042E3D3AD0C618B652A = I3C78D9AB59D6164851A819C5BA6C7C04 ;
assign I418D7ADEC09B065FFE6565D649D285B6 = IE12E3E0C53D89CE85C02DAFD3FB81244 ; assign IF2B42773D268BA706D29FCCFCB799AF9
= I8D8CDA8F60D3F8D5F51CD56B899536F8 ; assign I470C1C74A2768E559679EE12280C8506 = IC373345D0993637162B568673C9F7143 ;
assign I513461A4DA46CAA79BEC76A8DE8E2A98 = I5EBE440016CA0416EE3C2682065DDD85 ; assign ID7F4713F32DABD57E54222A946FA802F
= 1'b0; assign IADE62F3832E7DA9091E0F5B2EBC50F9C = 1'b0; assign I3443654006276E8DC7EE67AAE2283C64 = 1'b0; assign
I4FD27244D7DB92B0548A7AE35BDEDE28 = 1'b0; assign IDB44E9A441DC017FFA044AB8E232791F = (I569BD691A4BB295D836212F3738D46B4
== IE52A4905856745CF06589D8BBCBF62C0 ) ? 1'b1 : 1'b0;  assign ID59D28ABECF4E3544E08856EFCBC426D = I7EAA8AFFB2BC9D190B3626833AF5EBD8 ;
assign IE31D0AF3EFB3124913CD965CEE542B24 = IA21F6AD8A9BCF2140ECB6EE68E7A9FC5 & ~I928068FFB24833BA6A7A11BA59B8E040 ;
assign IA21F6AD8A9BCF2140ECB6EE68E7A9FC5 = (I3C78D9AB59D6164851A819C5BA6C7C04 == 2'b00) ? 1'b1 : ((I3C78D9AB59D6164851A819C5BA6C7C04
== 2'b01) ? I45917910AA4CC0F07BA1A8EF74FE6FEF [2] : I45917910AA4CC0F07BA1A8EF74FE6FEF [0]); assign I7EAA8AFFB2BC9D190B3626833AF5EBD8
= I06326CB6C7B31C2BC01AEF85D6548C61 | IADC13C79970748AA5DA1B07EC1C4290D | ICDFC5D4FA0C2CE90CDF9381D077D8CE2 | I756CF2AA8135461091FB5662DDE3111E ;
 always @(*) begin IFC499732997C1DCC89CB1F5E9F9C4CB3 = I569BD691A4BB295D836212F3738D46B4 ; case (I569BD691A4BB295D836212F3738D46B4 )
IC8B5868CE6CCCFF479B9D42AE258A6C9 : begin if (~I3E8F0524CDEE96F573376A6BF670184B ) IFC499732997C1DCC89CB1F5E9F9C4CB3
= IE52A4905856745CF06589D8BBCBF62C0 ; end IE52A4905856745CF06589D8BBCBF62C0 : begin IFC499732997C1DCC89CB1F5E9F9C4CB3
= I797FF78A781B011D1491E42DA6E8E636 ; end I797FF78A781B011D1491E42DA6E8E636 : begin if (I17066520A25539E7F98555DFF7832BBE
== 1'b1) IFC499732997C1DCC89CB1F5E9F9C4CB3 = I1829FA88EF5AD31D47831CE2250D10F7 ; end I1829FA88EF5AD31D47831CE2250D10F7
: begin IFC499732997C1DCC89CB1F5E9F9C4CB3 = IFCC4638207CC2B4943B7A3D236493B68 ; end IFCC4638207CC2B4943B7A3D236493B68
: begin if (I3565B787C28964F625269B34EE86A5CA ) IFC499732997C1DCC89CB1F5E9F9C4CB3 = I60218F936AC6C7F041F5C51CF271A588 ;
end I60218F936AC6C7F041F5C51CF271A588 : begin if (IABD5FBD9A9966396ACABECC997D287C6 & IFCFFF8448F5E6821B40C6CEE3548693A
& I7EAA8AFFB2BC9D190B3626833AF5EBD8 ) IFC499732997C1DCC89CB1F5E9F9C4CB3 = IB784FFF6C985E87492B9D6F18C3910AE ; end
IB784FFF6C985E87492B9D6F18C3910AE : begin if (IFCFFF8448F5E6821B40C6CEE3548693A ) if (I68014B0A38604EDB8B664C2C5CD25C03 )
IFC499732997C1DCC89CB1F5E9F9C4CB3 = I4ACB8367D46F2FB66718F5798E1F145F ; else IFC499732997C1DCC89CB1F5E9F9C4CB3 =
I293F67166A255C4EDC66C70F19551F8E ; end I293F67166A255C4EDC66C70F19551F8E : begin if (I68014B0A38604EDB8B664C2C5CD25C03
& IFCFFF8448F5E6821B40C6CEE3548693A ) IFC499732997C1DCC89CB1F5E9F9C4CB3 = I4ACB8367D46F2FB66718F5798E1F145F ; end
I4ACB8367D46F2FB66718F5798E1F145F : begin if (IFCFFF8448F5E6821B40C6CEE3548693A ) IFC499732997C1DCC89CB1F5E9F9C4CB3
= IC8B5868CE6CCCFF479B9D42AE258A6C9 ; end default : begin end endcase end  always @(*) begin case (I91A6742D4BEEA347CB6EDF3386EC70F6 )
I83EA49D19551ED8C672BF332D148F920 : begin IBC3E292376641E5290114F38B65B8702 = I2687BB96A4E1D15035B283D3FDF616CC ;
I68014B0A38604EDB8B664C2C5CD25C03 = IC4019EF7E804F3D95AAA442EFE259D86 ; end I373604D502FD927695BB13BAA1D3443F :
begin IBC3E292376641E5290114F38B65B8702 = I2EF8304B3AEA32E6C6F568223FAD9CBA ; I68014B0A38604EDB8B664C2C5CD25C03
= I8488C49C8D5977759183D4580A2BF116 ; end IA687834EBB97378F700DB12C9394F09F : begin IBC3E292376641E5290114F38B65B8702
= I369C6CA451B73B45E1F8D4D8AA53C2AD ; I68014B0A38604EDB8B664C2C5CD25C03 = I029FEAF1B2BC1E56CC9E23C77E352703 ; end
IF59ACE7A9B4E430EAAD83B6808CA927D : begin IBC3E292376641E5290114F38B65B8702 = IE81278F89BAA90C1F6EF0784D0DE2F62 ;
I68014B0A38604EDB8B664C2C5CD25C03 = IE4A11C65C530DD3B14BE1A05F3324401 ; end default : begin IBC3E292376641E5290114F38B65B8702
= {64{1'b0}}; I68014B0A38604EDB8B664C2C5CD25C03 = 1'b0; end endcase end  always @(posedge ICCFB0F435B37370076102F325BC08D20
or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin if (~I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin I31C96A05CDA83684954EE47D715D4665
<= 13'b0; I8E17DAB6BBC782E384ABBDDC296D791C <= 13'b0; I3565B787C28964F625269B34EE86A5CA <= 1'b0; IDA82F4C78A43B62E1C09ED19A1443221
<= 1'b0; IF4B2F356412545C21578876129150C2F <= 1'b0; I928068FFB24833BA6A7A11BA59B8E040 <= 1'b0; IE5C1CB646B621DD5D037AA5F5961D901
<= 64'b0; I1742675C5CD0344DCC6E13EC6252ED0A <= 1'b0; I23A5651CB59E99C9EF06BE735CE54321 <= 1'b0; IA1961DC2B849519BBCB37762269BB321
<= 1'b0; I9B1524315BD1F28EE8423E6A4D5CA375 <= 1'b0; I9A1E8CC9229E6A5D88D5CD96FBFE935D <= 1'b0; I637157BC0B4BC09421F86528FA1C6F22
<= 3'b0; I4DF8AE19A28761F0B98980365AEA794E <= 1'b0; I28BEA4229042F20DC4BAC5A80E0CF354 <= 10'b0; I6513C757AD9B98D491547EBB8D69BC7D
<= 1'b0; I297D3FE7B056FB743893BCFC1B67D805 <= 1'b0; I4F5985BF6243B7F0468BA4DD2B5D2E06 <= 1'b0; I3C78D9AB59D6164851A819C5BA6C7C04
<= 2'b00; IE12E3E0C53D89CE85C02DAFD3FB81244 <= 1'b0; I8D8CDA8F60D3F8D5F51CD56B899536F8 <= 1'b0; IC373345D0993637162B568673C9F7143
<= 1'b0; I5EBE440016CA0416EE3C2682065DDD85 <= 1'b0; IAA1E53CD0AE56DE019EFC1482B0134D6 <= 64'b0; I202B51CA022B3340D53544DEDC73872F
<= 64'b0; I37215D983C07F0C522E39A48B1F83101 <= 64'b0; I1F1327610E72511D7678CF70DE3685C6 <= 64'b0; I41D6A7D674F63A59E5DBBE00AA282E14
<= 1'b0; I23B9845BB3A093CE647D68158F400F36 <= 1'b0; I9542E55FC3D72D91960B79EC50367A55 <= 1'b0; I0CA51557A90D8B4060C406DC652C2485
<= 1'b0; I91A6742D4BEEA347CB6EDF3386EC70F6 <= 2'b0; I569BD691A4BB295D836212F3738D46B4 <= IC8B5868CE6CCCFF479B9D42AE258A6C9 ;
I45917910AA4CC0F07BA1A8EF74FE6FEF <= 3'b0; end else begin I31C96A05CDA83684954EE47D715D4665 <= I488999E90FEFB5E25518723EB6105532 ;
I8E17DAB6BBC782E384ABBDDC296D791C <= IA29842BA67669CD8D75483E633C363F0 ; I928068FFB24833BA6A7A11BA59B8E040 <= (IABD5FBD9A9966396ACABECC997D287C6
& IA21F6AD8A9BCF2140ECB6EE68E7A9FC5 ) | (I928068FFB24833BA6A7A11BA59B8E040 & ~(IFCFFF8448F5E6821B40C6CEE3548693A
& I23A5651CB59E99C9EF06BE735CE54321 )); I23A5651CB59E99C9EF06BE735CE54321 <= 1'b0; I9B1524315BD1F28EE8423E6A4D5CA375
<= 1'b0; I9A1E8CC9229E6A5D88D5CD96FBFE935D <= IFCFFF8448F5E6821B40C6CEE3548693A ; I637157BC0B4BC09421F86528FA1C6F22
<= I5CE5D2469FD5560C1773C754FC1E0C4A ; I4DF8AE19A28761F0B98980365AEA794E <= ID965E2D89D1047516134A3EED50CB8AE ;
IE12E3E0C53D89CE85C02DAFD3FB81244 <= 1'b0; I8D8CDA8F60D3F8D5F51CD56B899536F8 <= 1'b0; IC373345D0993637162B568673C9F7143
<= 1'b0; I5EBE440016CA0416EE3C2682065DDD85 <= 1'b0; IAA1E53CD0AE56DE019EFC1482B0134D6 <= I2687BB96A4E1D15035B283D3FDF616CC ;
I202B51CA022B3340D53544DEDC73872F <= I2EF8304B3AEA32E6C6F568223FAD9CBA ; I37215D983C07F0C522E39A48B1F83101 <= I369C6CA451B73B45E1F8D4D8AA53C2AD ;
I1F1327610E72511D7678CF70DE3685C6 <= IE81278F89BAA90C1F6EF0784D0DE2F62 ; I41D6A7D674F63A59E5DBBE00AA282E14 <= ~I2F86B5F8620848A51ED4F1F736CF8825 ;
I23B9845BB3A093CE647D68158F400F36 <= ~I63FDDFAA5AB093F3BB343A8C133F3BAF ; I9542E55FC3D72D91960B79EC50367A55 <= ~IE7F8A35B24BC8805CAD86FD378C18296 ;
I0CA51557A90D8B4060C406DC652C2485 <= ~IAB90D3559ED5004EBCCD9D73A2928E3F ; I6513C757AD9B98D491547EBB8D69BC7D <= (IAA1E53CD0AE56DE019EFC1482B0134D6 [1:0]
== 2'b0) ? ((I31C96A05CDA83684954EE47D715D4665 >= IAA1E53CD0AE56DE019EFC1482B0134D6 [9:2]) ? I41D6A7D674F63A59E5DBBE00AA282E14
: 1'b0) : ((I31C96A05CDA83684954EE47D715D4665 > IAA1E53CD0AE56DE019EFC1482B0134D6 [9:2]) ? I41D6A7D674F63A59E5DBBE00AA282E14
: 1'b0); I297D3FE7B056FB743893BCFC1B67D805 <= (I37215D983C07F0C522E39A48B1F83101 [1:0] == 2'b0) ? ((I8E17DAB6BBC782E384ABBDDC296D791C
>= I37215D983C07F0C522E39A48B1F83101 [9:2]) ? I9542E55FC3D72D91960B79EC50367A55 : 1'b0) : ((I8E17DAB6BBC782E384ABBDDC296D791C
> I37215D983C07F0C522E39A48B1F83101 [9:2]) ? I9542E55FC3D72D91960B79EC50367A55 : 1'b0); I4F5985BF6243B7F0468BA4DD2B5D2E06
<= (I1F1327610E72511D7678CF70DE3685C6 [1:0] == 2'b0) ? ((I8E17DAB6BBC782E384ABBDDC296D791C >= I1F1327610E72511D7678CF70DE3685C6 [9:2])
? I0CA51557A90D8B4060C406DC652C2485 : 1'b0) : ((I8E17DAB6BBC782E384ABBDDC296D791C > I1F1327610E72511D7678CF70DE3685C6 [9:2])
? I0CA51557A90D8B4060C406DC652C2485 : 1'b0); I45917910AA4CC0F07BA1A8EF74FE6FEF <= {I45917910AA4CC0F07BA1A8EF74FE6FEF [1:0],
IFCFFF8448F5E6821B40C6CEE3548693A }; I569BD691A4BB295D836212F3738D46B4 <= IFC499732997C1DCC89CB1F5E9F9C4CB3 ; if
(I4DF8AE19A28761F0B98980365AEA794E == 1'b0) case (I637157BC0B4BC09421F86528FA1C6F22 ) 3'b010 : I3C78D9AB59D6164851A819C5BA6C7C04
<= 2'b01; 3'b100 : I3C78D9AB59D6164851A819C5BA6C7C04 <= 2'b00; default : I3C78D9AB59D6164851A819C5BA6C7C04 <= 2'b10;
endcase else case (I637157BC0B4BC09421F86528FA1C6F22 ) 3'b010 : I3C78D9AB59D6164851A819C5BA6C7C04 <= 2'b00; default
: I3C78D9AB59D6164851A819C5BA6C7C04 <= 2'b01; endcase if (ID59D28ABECF4E3544E08856EFCBC426D == 1'b1) begin IE5C1CB646B621DD5D037AA5F5961D901
<= IBC3E292376641E5290114F38B65B8702 ; I1742675C5CD0344DCC6E13EC6252ED0A <= (I68014B0A38604EDB8B664C2C5CD25C03 ==
1'b0) ? 1'b0 : ((~IF4B2F356412545C21578876129150C2F & (~IDA82F4C78A43B62E1C09ED19A1443221 | ~I28BEA4229042F20DC4BAC5A80E0CF354 [0]))
| (IF4B2F356412545C21578876129150C2F & IDA82F4C78A43B62E1C09ED19A1443221 & I28BEA4229042F20DC4BAC5A80E0CF354 [0]));
end if (I17066520A25539E7F98555DFF7832BBE == 1'b1) I91A6742D4BEEA347CB6EDF3386EC70F6 <= I75EB9BE30F2D20C56659251E3B505209 ;
case (I569BD691A4BB295D836212F3738D46B4 ) IE52A4905856745CF06589D8BBCBF62C0 : begin I3565B787C28964F625269B34EE86A5CA
<= 1'b0; end I1829FA88EF5AD31D47831CE2250D10F7 : begin IDA82F4C78A43B62E1C09ED19A1443221 <= ((I91A6742D4BEEA347CB6EDF3386EC70F6
== I83EA49D19551ED8C672BF332D148F920 ) || (I91A6742D4BEEA347CB6EDF3386EC70F6 == IA687834EBB97378F700DB12C9394F09F )
|| (I91A6742D4BEEA347CB6EDF3386EC70F6 == IF59ACE7A9B4E430EAAD83B6808CA927D )) ? IBC3E292376641E5290114F38B65B8702 [62]
: 1'b0; IF4B2F356412545C21578876129150C2F <= ((I91A6742D4BEEA347CB6EDF3386EC70F6 == I373604D502FD927695BB13BAA1D3443F )
|| (I91A6742D4BEEA347CB6EDF3386EC70F6 == IA687834EBB97378F700DB12C9394F09F ) || (I91A6742D4BEEA347CB6EDF3386EC70F6
== IF59ACE7A9B4E430EAAD83B6808CA927D )) ? IBC3E292376641E5290114F38B65B8702 [61] : 1'b0; I28BEA4229042F20DC4BAC5A80E0CF354
<= IBC3E292376641E5290114F38B65B8702 [41:32]; end IFCC4638207CC2B4943B7A3D236493B68 : begin IA1961DC2B849519BBCB37762269BB321
<= I3565B787C28964F625269B34EE86A5CA ; case (I91A6742D4BEEA347CB6EDF3386EC70F6 ) I83EA49D19551ED8C672BF332D148F920
: begin if (IDA82F4C78A43B62E1C09ED19A1443221 ) I3565B787C28964F625269B34EE86A5CA <= (|IB064E00468F70C38840D1D271524C6C8 )
? I6513C757AD9B98D491547EBB8D69BC7D : 1'b0; else I3565B787C28964F625269B34EE86A5CA <= (|IB064E00468F70C38840D1D271524C6C8 )
? 1'b1 : 1'b0; end I373604D502FD927695BB13BAA1D3443F : begin I3565B787C28964F625269B34EE86A5CA <= (|I537C738B170D60A42A1F6FDA4547BACC )
? 1'b1 : 1'b0; end IA687834EBB97378F700DB12C9394F09F : begin if (IDA82F4C78A43B62E1C09ED19A1443221 ) I3565B787C28964F625269B34EE86A5CA
<= (|IB9E3BDBEE7C442BA69CD12711DA40F71 ) ? I297D3FE7B056FB743893BCFC1B67D805 : 1'b0; else I3565B787C28964F625269B34EE86A5CA
<= (|IB9E3BDBEE7C442BA69CD12711DA40F71 ) ? 1'b1 : 1'b0; end IF59ACE7A9B4E430EAAD83B6808CA927D : begin if (IDA82F4C78A43B62E1C09ED19A1443221 )
I3565B787C28964F625269B34EE86A5CA <= (|IB9E3BDBEE7C442BA69CD12711DA40F71 ) ? I4F5985BF6243B7F0468BA4DD2B5D2E06 :
1'b0; else I3565B787C28964F625269B34EE86A5CA <= (|IB9E3BDBEE7C442BA69CD12711DA40F71 ) ? 1'b1 : 1'b0; end endcase
end I60218F936AC6C7F041F5C51CF271A588 : begin IA1961DC2B849519BBCB37762269BB321 <= IA1961DC2B849519BBCB37762269BB321
& ~(IABD5FBD9A9966396ACABECC997D287C6 & IFCFFF8448F5E6821B40C6CEE3548693A ); I9B1524315BD1F28EE8423E6A4D5CA375 <=
I7EAA8AFFB2BC9D190B3626833AF5EBD8 ;   IE12E3E0C53D89CE85C02DAFD3FB81244 <= (I91A6742D4BEEA347CB6EDF3386EC70F6 ==
I83EA49D19551ED8C672BF332D148F920 ) ? (IABD5FBD9A9966396ACABECC997D287C6 & IE31D0AF3EFB3124913CD965CEE542B24 ) :
1'b0; I8D8CDA8F60D3F8D5F51CD56B899536F8 <= (I91A6742D4BEEA347CB6EDF3386EC70F6 == I373604D502FD927695BB13BAA1D3443F )
? (IABD5FBD9A9966396ACABECC997D287C6 & IE31D0AF3EFB3124913CD965CEE542B24 ) : 1'b0; IC373345D0993637162B568673C9F7143
<= (I91A6742D4BEEA347CB6EDF3386EC70F6 == IA687834EBB97378F700DB12C9394F09F ) ? (IABD5FBD9A9966396ACABECC997D287C6
& IE31D0AF3EFB3124913CD965CEE542B24 ) : 1'b0; I5EBE440016CA0416EE3C2682065DDD85 <= (I91A6742D4BEEA347CB6EDF3386EC70F6
== IF59ACE7A9B4E430EAAD83B6808CA927D ) ? (IABD5FBD9A9966396ACABECC997D287C6 & IE31D0AF3EFB3124913CD965CEE542B24 )
: 1'b0; end IB784FFF6C985E87492B9D6F18C3910AE : begin I23A5651CB59E99C9EF06BE735CE54321 <= I68014B0A38604EDB8B664C2C5CD25C03
& IFCFFF8448F5E6821B40C6CEE3548693A ; I9B1524315BD1F28EE8423E6A4D5CA375 <= I9B1524315BD1F28EE8423E6A4D5CA375 & ~IFCFFF8448F5E6821B40C6CEE3548693A ;
end I293F67166A255C4EDC66C70F19551F8E : begin I23A5651CB59E99C9EF06BE735CE54321 <= I68014B0A38604EDB8B664C2C5CD25C03
& IFCFFF8448F5E6821B40C6CEE3548693A ; end I4ACB8367D46F2FB66718F5798E1F145F : begin I23A5651CB59E99C9EF06BE735CE54321
<= I23A5651CB59E99C9EF06BE735CE54321 & ~IFCFFF8448F5E6821B40C6CEE3548693A ; end endcase end end endmodule 
  module I1D0F7B4B91A0FA84F3F3816624A1A70F #( parameter I87C69AEB153025D890F0A7CE399F00FE = 3 ) ( input wire ICCFB0F435B37370076102F325BC08D20 ,
input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire IBA6CF56719009F0FF759C0AF1F1630AF , input wire I42D2723FE4CDE4AF565DD01BD32BB8AC ,
input wire I8E99DEF5C63C6A55606BD30E4BE8E3FB , input wire IC3760F6E74F9AA61561390CC1466FC1A , input wire I582940C94DBA710A62923187D833E8E6 ,
output wire IAFF3235BDF22DE6B7D7DBF12451FA2FE , output wire I5FFD1878342C11E50C1617928EBB38D7 , output wire I27766E6DFBDE7E37CDB16F4E2C0E1DD4 ,
output wire I520751EAD225B5BFC3D7E0ACB7BC6405 , output wire [I87C69AEB153025D890F0A7CE399F00FE - 1:0] I94ED0A1B920B23A4D17502C81A2A18C7 ,
output wire I6010C20131B976554A498745FEEEB580 ); `include "tlp_qcodes.v"
 reg I29050B07476020B7A718339867806908 ; reg IFC73E93AA35A80792ADE9017768129C1 ; reg I525B2ED0A58FC2F85C15158BA3F67357 ;
reg I48F84F9DB41F3E71C472A13B0AD06720 ; reg I5B3BB6CF473F793585E2668A9A7136C8 ; reg [I87C69AEB153025D890F0A7CE399F00FE
- 1:0] IBE3F740634E17CD7B70D2C7ACCB20B8F ; wire [3:0] IDD1B0C54E1662B5BFB789B4A625CECAD ;  assign IAFF3235BDF22DE6B7D7DBF12451FA2FE
= I29050B07476020B7A718339867806908 ; assign I5FFD1878342C11E50C1617928EBB38D7 = IFC73E93AA35A80792ADE9017768129C1 ;
assign I27766E6DFBDE7E37CDB16F4E2C0E1DD4 = I525B2ED0A58FC2F85C15158BA3F67357 ; assign I520751EAD225B5BFC3D7E0ACB7BC6405
= I48F84F9DB41F3E71C472A13B0AD06720 ; assign I6010C20131B976554A498745FEEEB580 = I5B3BB6CF473F793585E2668A9A7136C8 ;
assign I94ED0A1B920B23A4D17502C81A2A18C7 = IBE3F740634E17CD7B70D2C7ACCB20B8F ;   assign IDD1B0C54E1662B5BFB789B4A625CECAD
= {I8E99DEF5C63C6A55606BD30E4BE8E3FB , I582940C94DBA710A62923187D833E8E6 , I42D2723FE4CDE4AF565DD01BD32BB8AC , IC3760F6E74F9AA61561390CC1466FC1A };
 always @(posedge ICCFB0F435B37370076102F325BC08D20 or negedge I9ED2A9117D3AEAF54CBA7AD69083BCB7 ) begin if (~I9ED2A9117D3AEAF54CBA7AD69083BCB7 )
begin I29050B07476020B7A718339867806908 <= 1'b0; IFC73E93AA35A80792ADE9017768129C1 <= 1'b0; I525B2ED0A58FC2F85C15158BA3F67357
<= 1'b0; I48F84F9DB41F3E71C472A13B0AD06720 <= 1'b0; I5B3BB6CF473F793585E2668A9A7136C8 <= 1'b0; IBE3F740634E17CD7B70D2C7ACCB20B8F
<= {I87C69AEB153025D890F0A7CE399F00FE {1'b0}}; end else begin I29050B07476020B7A718339867806908 <= 1'b0; IFC73E93AA35A80792ADE9017768129C1
<= 1'b0; I525B2ED0A58FC2F85C15158BA3F67357 <= 1'b0; I48F84F9DB41F3E71C472A13B0AD06720 <= 1'b0; I5B3BB6CF473F793585E2668A9A7136C8
<= 1'b0; IBE3F740634E17CD7B70D2C7ACCB20B8F <= {I87C69AEB153025D890F0A7CE399F00FE {1'b0}}; casex (IDD1B0C54E1662B5BFB789B4A625CECAD )
4'bxxx1 : begin I525B2ED0A58FC2F85C15158BA3F67357 <= IC3760F6E74F9AA61561390CC1466FC1A & ~(IBA6CF56719009F0FF759C0AF1F1630AF
| I5B3BB6CF473F793585E2668A9A7136C8 ); I5B3BB6CF473F793585E2668A9A7136C8 <= ~(IBA6CF56719009F0FF759C0AF1F1630AF
| I5B3BB6CF473F793585E2668A9A7136C8 ); IBE3F740634E17CD7B70D2C7ACCB20B8F <= IA687834EBB97378F700DB12C9394F09F ;
end 4'bxx10 : begin I29050B07476020B7A718339867806908 <= I42D2723FE4CDE4AF565DD01BD32BB8AC & ~(IBA6CF56719009F0FF759C0AF1F1630AF
| I5B3BB6CF473F793585E2668A9A7136C8 ); I5B3BB6CF473F793585E2668A9A7136C8 <= ~(IBA6CF56719009F0FF759C0AF1F1630AF
| I5B3BB6CF473F793585E2668A9A7136C8 ); IBE3F740634E17CD7B70D2C7ACCB20B8F <= I83EA49D19551ED8C672BF332D148F920 ;
end 4'bx100 : begin I48F84F9DB41F3E71C472A13B0AD06720 <= I582940C94DBA710A62923187D833E8E6 & ~(IBA6CF56719009F0FF759C0AF1F1630AF
| I5B3BB6CF473F793585E2668A9A7136C8 ); I5B3BB6CF473F793585E2668A9A7136C8 <= ~(IBA6CF56719009F0FF759C0AF1F1630AF
| I5B3BB6CF473F793585E2668A9A7136C8 ); IBE3F740634E17CD7B70D2C7ACCB20B8F <= IF59ACE7A9B4E430EAAD83B6808CA927D ;
end 4'b1000 : begin IFC73E93AA35A80792ADE9017768129C1 <= I8E99DEF5C63C6A55606BD30E4BE8E3FB & ~(IBA6CF56719009F0FF759C0AF1F1630AF
| I5B3BB6CF473F793585E2668A9A7136C8 ); I5B3BB6CF473F793585E2668A9A7136C8 <= ~(IBA6CF56719009F0FF759C0AF1F1630AF
| I5B3BB6CF473F793585E2668A9A7136C8 ); IBE3F740634E17CD7B70D2C7ACCB20B8F <= I373604D502FD927695BB13BAA1D3443F ;
end default : begin end endcase end end endmodule
  module ICF327C89C36124513E146F1FF3BCDEEB #( parameter I87C69AEB153025D890F0A7CE399F00FE = 3, parameter I68B4790A0165FFB6E2740B409126FE6B
= 8, I66C185998F46A7148163982E39BCD296 = "ecp3" )( input wire ICCFB0F435B37370076102F325BC08D20 , input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 ,
input wire I0C5BEBB297319D36CFD96B791AFE888C , input wire I42D2723FE4CDE4AF565DD01BD32BB8AC , input wire I8E99DEF5C63C6A55606BD30E4BE8E3FB ,
input wire IC3760F6E74F9AA61561390CC1466FC1A , input wire I582940C94DBA710A62923187D833E8E6 , output wire IAFF3235BDF22DE6B7D7DBF12451FA2FE ,
output wire I5FFD1878342C11E50C1617928EBB38D7 , output wire I27766E6DFBDE7E37CDB16F4E2C0E1DD4 , output wire I520751EAD225B5BFC3D7E0ACB7BC6405 ,
output wire [I87C69AEB153025D890F0A7CE399F00FE - 1:0] IFA5857E29877E868702F9890224BA5FC , output wire I3CEE775C269D38D2B516507E40A6387C ,
output wire IEADE52DA6BAC6B55AC606944635D8C9A );  wire IA83F679A674E1F4A4A69FDB86C6E339F ; wire I5564F0E4F9AE04792C7CCADA977449AD ;
wire I932E68CEB931A44CEF843351FD7AA7D0 ; wire IFED7584192506445FFD17C3921381807 ; wire I4DDC35D2ABD8CA6BE29CAC68BC10C340 ;
wire [I87C69AEB153025D890F0A7CE399F00FE - 1:0] ID20B34301F6953CD6F5008CB3B6A369A ; wire [I87C69AEB153025D890F0A7CE399F00FE
- 1:0] I45B614E1199C70B4E5F58D3EFD1D08C7 ; wire I69B84382CF4434D3BBB964B953CD6E15 ; wire IE24F5745323EB576C5BF2A24254B882B ;
wire IE61B38939030FBBD451B170FB1F376E7 ;  assign IAFF3235BDF22DE6B7D7DBF12451FA2FE = IA83F679A674E1F4A4A69FDB86C6E339F ;
assign I5FFD1878342C11E50C1617928EBB38D7 = I5564F0E4F9AE04792C7CCADA977449AD ; assign I27766E6DFBDE7E37CDB16F4E2C0E1DD4
= I932E68CEB931A44CEF843351FD7AA7D0 ; assign I520751EAD225B5BFC3D7E0ACB7BC6405 = IFED7584192506445FFD17C3921381807 ;
assign IFA5857E29877E868702F9890224BA5FC = I45B614E1199C70B4E5F58D3EFD1D08C7 ; assign I3CEE775C269D38D2B516507E40A6387C
= I69B84382CF4434D3BBB964B953CD6E15 ; assign IEADE52DA6BAC6B55AC606944635D8C9A = IE61B38939030FBBD451B170FB1F376E7 ;
 I1D0F7B4B91A0FA84F3F3816624A1A70F #( .I87C69AEB153025D890F0A7CE399F00FE (I87C69AEB153025D890F0A7CE399F00FE ) )
IB420C4D1279F971E867FA537CA4D6E82 ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .IBA6CF56719009F0FF759C0AF1F1630AF (IE24F5745323EB576C5BF2A24254B882B ), .I42D2723FE4CDE4AF565DD01BD32BB8AC
(I42D2723FE4CDE4AF565DD01BD32BB8AC ), .I8E99DEF5C63C6A55606BD30E4BE8E3FB (I8E99DEF5C63C6A55606BD30E4BE8E3FB ), .IC3760F6E74F9AA61561390CC1466FC1A
(IC3760F6E74F9AA61561390CC1466FC1A ), .I582940C94DBA710A62923187D833E8E6 (I582940C94DBA710A62923187D833E8E6 ), .IAFF3235BDF22DE6B7D7DBF12451FA2FE
(IA83F679A674E1F4A4A69FDB86C6E339F ), .I5FFD1878342C11E50C1617928EBB38D7 (I5564F0E4F9AE04792C7CCADA977449AD ), .I27766E6DFBDE7E37CDB16F4E2C0E1DD4
(I932E68CEB931A44CEF843351FD7AA7D0 ), .I520751EAD225B5BFC3D7E0ACB7BC6405 (IFED7584192506445FFD17C3921381807 ), .I94ED0A1B920B23A4D17502C81A2A18C7
(ID20B34301F6953CD6F5008CB3B6A369A ), .I6010C20131B976554A498745FEEEB580 (I4DDC35D2ABD8CA6BE29CAC68BC10C340 ) );
IF4FD65273243DC47A72869EEEA639DCD #( .I7292F55C07BFD7FB8A60D29FFC186275 (I87C69AEB153025D890F0A7CE399F00FE ), .IB71844FFA3AB85FEF45EAB4D35395752
(I68B4790A0165FFB6E2740B409126FE6B ), .I66C185998F46A7148163982E39BCD296 (I66C185998F46A7148163982E39BCD296 ) )
IA440041682C400211AAD0D987978451E ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .IC79EC9A9F373F4B71374BDF6EDD31DE6 (1'b0), .I48D61F5A0B5732A58912433B42CD9D0C
(I0C5BEBB297319D36CFD96B791AFE888C ), .I04BC24D2B6403E54A64DE9E6C9ABAA2B (ID20B34301F6953CD6F5008CB3B6A369A ), .IE315CDCA06C9620D5C0AB966E553F0C3
(I4DDC35D2ABD8CA6BE29CAC68BC10C340 ), .I11CEFC90537A67CD1FF01400245362F2 ( ), .ID7FCE45A65ADDB17F91F73A1B506BB5B
( ), .I125028C7446331521D0434C10E8B0007 (I45B614E1199C70B4E5F58D3EFD1D08C7 ), .I8BB939FF2AFDE7B2A1E480DCB61CE354
(I69B84382CF4434D3BBB964B953CD6E15 ), .I41C63F948E534C7ED9F2471A44C922B2 ( ), .I585F74DE05DD9C1C7070D6B4F6E181C2
(IE61B38939030FBBD451B170FB1F376E7 ), .I705C64753A50CDA034B5ACB332D71768 ( ), .I233E0C0C8E5150F0CD8258F276D93942
( ), .IBE0D6810EBD63B5C428623C578CF6D3A (IE24F5745323EB576C5BF2A24254B882B ), .I115E90220158F08B0465E99D7F2561D3
( ) ); endmodule 
  `timescale 1 ns / 1 ps 
module I7639B3DE6448BF04A6DF404C0FEDBA75 #( parameter I7292F55C07BFD7FB8A60D29FFC186275 = 32, parameter IDB751C3DD512B8355CF27001F983880A
= 16, parameter I99651B9F47529E0ADC5349B57C84E531 = 512, parameter ICED1C5B792370B25488CFA18FE5E472E = 512, parameter
I0AEF008AE3BC7E23C49F86BC2B344750 = 512, parameter I026FA76AB836F95856A0F400EDF284FA = 512, parameter I66C185998F46A7148163982E39BCD296
= "ecp3", parameter I6684631E4DAAC3FB7551EF267A7E3D73 = 32, parameter I3A59A966031A54015DBF77A68A5A82D3 = 32 ) (
input wire ICCFB0F435B37370076102F325BC08D20 , input wire I9ED2A9117D3AEAF54CBA7AD69083BCB7 , input wire [12:0]
I488999E90FEFB5E25518723EB6105532 , input wire [8:0] IB064E00468F70C38840D1D271524C6C8 , input wire [12:0] IE4E19EA6F3F828B3B44ED1E4D36558F7 ,
input wire [8:0] I537C738B170D60A42A1F6FDA4547BACC , input wire [12:0] IA29842BA67669CD8D75483E633C363F0 , input
wire [8:0] IB9E3BDBEE7C442BA69CD12711DA40F71 , input wire IABD5FBD9A9966396ACABECC997D287C6 , input wire IFCFFF8448F5E6821B40C6CEE3548693A ,
input wire [2:0] I5CE5D2469FD5560C1773C754FC1E0C4A , input wire ID965E2D89D1047516134A3EED50CB8AE , input wire [I6684631E4DAAC3FB7551EF267A7E3D73
- 1:0] I884F4ADE09FABBA20600F67BC1A50FE7 , input wire I61E8E6981294A3342BDF5596043A2DFA , input wire I2F5C52C0CABA5EFAF34A96BC39DA8F96 ,
input wire [I3A59A966031A54015DBF77A68A5A82D3 - 1:0] I0BA940AC86B853EFCE63667C128E2DF4 , input wire ID176017A6F96653AFD707B70D22BEA8C ,
input wire IE8C34BE7792A66A23CB1C7A5CFF55BBF , input wire [I6684631E4DAAC3FB7551EF267A7E3D73 - 1:0] IA5896E672427191F9A0B4ED1C9301313 ,
input wire I0317313DEECD8AC19E98BA2F1C27E0A9 , input wire IFDB2ACAC637F40CDDFBB20A3AFD9A401 , input wire [I3A59A966031A54015DBF77A68A5A82D3
- 1:0] IE4C3654339F6BF285840C2AB868371A1 , input wire I5F40D6DD3270B21E2E90925F127E6477 , input wire I33A8C146E90D24E54E605500849CD461 ,
input wire I42D2723FE4CDE4AF565DD01BD32BB8AC , input wire I8E99DEF5C63C6A55606BD30E4BE8E3FB , input wire IC3760F6E74F9AA61561390CC1466FC1A ,
input wire I582940C94DBA710A62923187D833E8E6 , output wire [$clog2((I99651B9F47529E0ADC5349B57C84E531 * (I7292F55C07BFD7FB8A60D29FFC186275 /I6684631E4DAAC3FB7551EF267A7E3D73 ))
+ 1) - 1:0] IDFCF1C6E3889548A5224E9568D7E2E22 , output wire [$clog2((ICED1C5B792370B25488CFA18FE5E472E * (I7292F55C07BFD7FB8A60D29FFC186275 /I6684631E4DAAC3FB7551EF267A7E3D73 ))
+ 1) - 1 : 0] I241490D6913C41E3972F651398E36880 , output wire [$clog2((I0AEF008AE3BC7E23C49F86BC2B344750 * (I7292F55C07BFD7FB8A60D29FFC186275 /I6684631E4DAAC3FB7551EF267A7E3D73 ))
+ 1) - 1 : 0] IA127FE276B1C05C6A690F8454BBF510B , output wire [$clog2((I026FA76AB836F95856A0F400EDF284FA * (I7292F55C07BFD7FB8A60D29FFC186275 /I6684631E4DAAC3FB7551EF267A7E3D73 ))
+ 1) - 1:0] I0ED116F3061ADCE682AE68F0A5003CBF , output wire [IDB751C3DD512B8355CF27001F983880A - 1:0] IB33B8D629A269D1BC3D79902EE2EB312 ,
output wire I1E494BBA2ECB063404DBB73667CC7E8D , output wire I4A4976CAF016EA789DCDB7AA131246C3 , output wire I5ADFC7E7F8B570F5258C2813D0020950 ,
output wire I1FD27F5D298FA5493F3F510610F19E4E , output wire IAFF3235BDF22DE6B7D7DBF12451FA2FE , output wire I5FFD1878342C11E50C1617928EBB38D7 ,
output wire I27766E6DFBDE7E37CDB16F4E2C0E1DD4 , output wire I520751EAD225B5BFC3D7E0ACB7BC6405 ); `include "tlp_qcodes.v"
 localparam I9C4BDAB65913DE43240C2A937C25DD0D = $clog2((I99651B9F47529E0ADC5349B57C84E531 * (I7292F55C07BFD7FB8A60D29FFC186275 /I6684631E4DAAC3FB7551EF267A7E3D73 ))
+ 1); localparam ICEFA062966B07CA76E008210CF0F32DC = $clog2((ICED1C5B792370B25488CFA18FE5E472E * (I7292F55C07BFD7FB8A60D29FFC186275 /I3A59A966031A54015DBF77A68A5A82D3 ))
+ 1); localparam IE823348F0219A94EDEF99E63176786C4 = $clog2((I0AEF008AE3BC7E23C49F86BC2B344750 * (I7292F55C07BFD7FB8A60D29FFC186275 /I6684631E4DAAC3FB7551EF267A7E3D73 ))
+ 1); localparam I96F78D1E32AB1DCE01DB91736CB0459C = $clog2((I026FA76AB836F95856A0F400EDF284FA * (I7292F55C07BFD7FB8A60D29FFC186275 /I3A59A966031A54015DBF77A68A5A82D3 ))
+ 1);  wire [IDB751C3DD512B8355CF27001F983880A - 1:0] IA69B6A69D96E898639A555BF6567C273 ; wire IFD8A5AA76F99D6914AE0274FCD000AD1 ;
wire ICA6FC4E4455EED217775291436AD860C ; wire IFE46A9371C863D1229E8DCA840188E17 ; wire IF63E39473014C2B5C4FB8832104F3754 ;
wire [1:0] I58FB5703785F6B602E564F2C3886577D ; wire IC85FD97ECAC87466B9C19ACECC79FC2D ; wire IA5B538B804B78BFE2529013B5C97D493 ;
wire IB7543BE04BDCE5E5193E442BACB25B09 ; wire IC6D81493F78B34E8262D34CE51650B27 ; wire ID40108F42D0FA32BFA839EFAD8F8C320 ;
wire I46618BF7FF1CE70399E81FFAD2D6846B ; wire I1CA27197DF7539251654AB3DAC8E8B38 ; wire I755156D55303F238FD088C21A8C23864 ;
wire ID2C4F123A6A9197C7B4B4FD780FCC272 ; wire I48ABEC51DF27ACA5596235F4DF0D08C4 ; wire IF77AAC35DEF2E12949B516C97BABF4FD ;
wire I586E9AE745283DB69A128B0C7A472DE0 ; wire I91383F42CED2732A542098CD5ACFFD1D ; wire [IC7701945BBBE654661A8C2F153881F63 :0]
I45B614E1199C70B4E5F58D3EFD1D08C7 ; wire I69B84382CF4434D3BBB964B953CD6E15 ; wire IF66089F4B958743DD8052C5F9D832CD1 ;
wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] I2F2159E4520CF0D6E57382C8E60EC46D ; wire I4DDF7CB99428D62C1FB17E5C8FA42E6A ;
wire [I9C4BDAB65913DE43240C2A937C25DD0D - 1:0] I7F72A1B5D33702E3B645BD20CB425937 ; wire IA4EA76535E7026B1F7DF3EDC236AF756 ;
wire I7DA036F5B0B44A1D5E3EB0237828A810 ; wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] I673AF3DF8D93FAFCF8E255C8C6852D9B ;
wire IB76DC52DFFF4905395FBC5C33F2C6B24 ; wire [IE823348F0219A94EDEF99E63176786C4 - 1:0] IB6FE1681C40869E515EA3BF2BD5F7DA8 ;
wire I9D0CEC2083A8932FA283AD091303049F ; wire IE43DA634E45C0D88369455568042AF37 ; wire [I7292F55C07BFD7FB8A60D29FFC186275
- 1:0] I2BE5B3BCC47A675D856661ED2CA18C19 ; wire I8236407E542CBF20A06054E415DF3019 ; wire [I96F78D1E32AB1DCE01DB91736CB0459C
- 1:0] I96EC08C26A305FC6029163D693EF44E6 ; wire I173FA018899178893FB946275729ED68 ; wire I5871F7D82773EB9D3EE955FCC1611D9F ;
wire [I7292F55C07BFD7FB8A60D29FFC186275 - 1:0] IC1C88613A52A238F417438A678D1196A ; wire I7B40A3A5ECAB9C16D0C5E2614F94A037 ;
wire [ICEFA062966B07CA76E008210CF0F32DC - 1:0] I5E12F1044C6612C74B661A7400A97D4B ; wire ID505752183B05B70B86F1045E7DB0CF0 ;
wire I36AD11753E1A0E22546912955186E616 ;  assign IDFCF1C6E3889548A5224E9568D7E2E22 = I7F72A1B5D33702E3B645BD20CB425937 ;
assign I241490D6913C41E3972F651398E36880 = I5E12F1044C6612C74B661A7400A97D4B ; assign IA127FE276B1C05C6A690F8454BBF510B
= IB6FE1681C40869E515EA3BF2BD5F7DA8 ; assign I0ED116F3061ADCE682AE68F0A5003CBF = I96EC08C26A305FC6029163D693EF44E6 ;
assign IB33B8D629A269D1BC3D79902EE2EB312 = IA69B6A69D96E898639A555BF6567C273 ; assign I1E494BBA2ECB063404DBB73667CC7E8D
= (IDB751C3DD512B8355CF27001F983880A == 16) ? 1'b0 : IFD8A5AA76F99D6914AE0274FCD000AD1 ; assign I4A4976CAF016EA789DCDB7AA131246C3
= ICA6FC4E4455EED217775291436AD860C ; assign I5ADFC7E7F8B570F5258C2813D0020950 = IFE46A9371C863D1229E8DCA840188E17 ;
assign I1FD27F5D298FA5493F3F510610F19E4E = IF63E39473014C2B5C4FB8832104F3754 ; assign IAFF3235BDF22DE6B7D7DBF12451FA2FE
= I48ABEC51DF27ACA5596235F4DF0D08C4 ; assign I5FFD1878342C11E50C1617928EBB38D7 = IF77AAC35DEF2E12949B516C97BABF4FD ;
assign I27766E6DFBDE7E37CDB16F4E2C0E1DD4 = I586E9AE745283DB69A128B0C7A472DE0 ; assign I520751EAD225B5BFC3D7E0ACB7BC6405
= I91383F42CED2732A542098CD5ACFFD1D ;  generate if (IDB751C3DD512B8355CF27001F983880A == 16) begin : IBC503D04A72C6E62ECAE6A99BC68A860
I8489B3291801D4F3BE8AED05E26C4566 #( .I87C69AEB153025D890F0A7CE399F00FE (IBACE8243A55E1A6C355E86BA25034EFB ) ) I052230D66B4BFAAC87011F404C4761F3
( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ),
.I488999E90FEFB5E25518723EB6105532 (I488999E90FEFB5E25518723EB6105532 ), .IB064E00468F70C38840D1D271524C6C8 (IB064E00468F70C38840D1D271524C6C8 ),
.IE4E19EA6F3F828B3B44ED1E4D36558F7 (IE4E19EA6F3F828B3B44ED1E4D36558F7 ), .I537C738B170D60A42A1F6FDA4547BACC (I537C738B170D60A42A1F6FDA4547BACC ),
.IA29842BA67669CD8D75483E633C363F0 (IA29842BA67669CD8D75483E633C363F0 ), .IB9E3BDBEE7C442BA69CD12711DA40F71 (IB9E3BDBEE7C442BA69CD12711DA40F71 ),
.IABD5FBD9A9966396ACABECC997D287C6 (IABD5FBD9A9966396ACABECC997D287C6 ), .I06326CB6C7B31C2BC01AEF85D6548C61 (I7DA036F5B0B44A1D5E3EB0237828A810 ),
.IADC13C79970748AA5DA1B07EC1C4290D (IE43DA634E45C0D88369455568042AF37 ), .ICDFC5D4FA0C2CE90CDF9381D077D8CE2 (I5871F7D82773EB9D3EE955FCC1611D9F ),
.I756CF2AA8135461091FB5662DDE3111E (I36AD11753E1A0E22546912955186E616 ), .I2687BB96A4E1D15035B283D3FDF616CC (I2F2159E4520CF0D6E57382C8E60EC46D ),
.I2EF8304B3AEA32E6C6F568223FAD9CBA (IC1C88613A52A238F417438A678D1196A ), .I369C6CA451B73B45E1F8D4D8AA53C2AD (I673AF3DF8D93FAFCF8E255C8C6852D9B ),
.IE81278F89BAA90C1F6EF0784D0DE2F62 (I2BE5B3BCC47A675D856661ED2CA18C19 ), .I2F86B5F8620848A51ED4F1F736CF8825 (I4DDF7CB99428D62C1FB17E5C8FA42E6A ),
.I63FDDFAA5AB093F3BB343A8C133F3BAF (I7B40A3A5ECAB9C16D0C5E2614F94A037 ), .IE7F8A35B24BC8805CAD86FD378C18296 (IB76DC52DFFF4905395FBC5C33F2C6B24 ),
.IAB90D3559ED5004EBCCD9D73A2928E3F (I8236407E542CBF20A06054E415DF3019 ), .I75EB9BE30F2D20C56659251E3B505209 (I45B614E1199C70B4E5F58D3EFD1D08C7 ),
.I3E8F0524CDEE96F573376A6BF670184B (I69B84382CF4434D3BBB964B953CD6E15 ), .I17066520A25539E7F98555DFF7832BBE (IF66089F4B958743DD8052C5F9D832CD1 ),
.IB33B8D629A269D1BC3D79902EE2EB312 (IA69B6A69D96E898639A555BF6567C273 ), .I4A4976CAF016EA789DCDB7AA131246C3 (ICA6FC4E4455EED217775291436AD860C ),
.I5ADFC7E7F8B570F5258C2813D0020950 (IFE46A9371C863D1229E8DCA840188E17 ), .I1FD27F5D298FA5493F3F510610F19E4E (IF63E39473014C2B5C4FB8832104F3754 ),
.ID7F4713F32DABD57E54222A946FA802F (ID40108F42D0FA32BFA839EFAD8F8C320 ), .IADE62F3832E7DA9091E0F5B2EBC50F9C (I46618BF7FF1CE70399E81FFAD2D6846B ),
.I3443654006276E8DC7EE67AAE2283C64 (I1CA27197DF7539251654AB3DAC8E8B38 ), .I4FD27244D7DB92B0548A7AE35BDEDE28 (I755156D55303F238FD088C21A8C23864 ),
.IDB44E9A441DC017FFA044AB8E232791F (ID2C4F123A6A9197C7B4B4FD780FCC272 ) ); assign IC85FD97ECAC87466B9C19ACECC79FC2D
= 1'b0; assign IB7543BE04BDCE5E5193E442BACB25B09 = 1'b0; assign IC6D81493F78B34E8262D34CE51650B27 = 1'b0; assign
IA5B538B804B78BFE2529013B5C97D493 = 1'b0; end endgenerate generate if (IDB751C3DD512B8355CF27001F983880A == 64)
begin : I9DEBD354280DD846EE864EC5E3157726 I5AA57FA362D8C2F14DF19B01C99AE372 #( .I87C69AEB153025D890F0A7CE399F00FE
(IBACE8243A55E1A6C355E86BA25034EFB ) ) I052230D66B4BFAAC87011F404C4761F3 ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ),
.I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .I488999E90FEFB5E25518723EB6105532 (I488999E90FEFB5E25518723EB6105532 ),
.IB064E00468F70C38840D1D271524C6C8 (IB064E00468F70C38840D1D271524C6C8 ), .IE4E19EA6F3F828B3B44ED1E4D36558F7 (IE4E19EA6F3F828B3B44ED1E4D36558F7 ),
.I537C738B170D60A42A1F6FDA4547BACC (I537C738B170D60A42A1F6FDA4547BACC ), .IA29842BA67669CD8D75483E633C363F0 (IA29842BA67669CD8D75483E633C363F0 ),
.IB9E3BDBEE7C442BA69CD12711DA40F71 (IB9E3BDBEE7C442BA69CD12711DA40F71 ), .IABD5FBD9A9966396ACABECC997D287C6 (IABD5FBD9A9966396ACABECC997D287C6 ),
.IFCFFF8448F5E6821B40C6CEE3548693A (IFCFFF8448F5E6821B40C6CEE3548693A ), .I5CE5D2469FD5560C1773C754FC1E0C4A (I5CE5D2469FD5560C1773C754FC1E0C4A ),
.ID965E2D89D1047516134A3EED50CB8AE (ID965E2D89D1047516134A3EED50CB8AE ), .IC4019EF7E804F3D95AAA442EFE259D86 (IA4EA76535E7026B1F7DF3EDC236AF756 ),
.I8488C49C8D5977759183D4580A2BF116 (ID505752183B05B70B86F1045E7DB0CF0 ), .I029FEAF1B2BC1E56CC9E23C77E352703 (I9D0CEC2083A8932FA283AD091303049F ),
.IE4A11C65C530DD3B14BE1A05F3324401 (I173FA018899178893FB946275729ED68 ), .I06326CB6C7B31C2BC01AEF85D6548C61 (I7DA036F5B0B44A1D5E3EB0237828A810 ),
.IADC13C79970748AA5DA1B07EC1C4290D (I36AD11753E1A0E22546912955186E616 ), .ICDFC5D4FA0C2CE90CDF9381D077D8CE2 (IE43DA634E45C0D88369455568042AF37 ),
.I756CF2AA8135461091FB5662DDE3111E (I5871F7D82773EB9D3EE955FCC1611D9F ), .I2687BB96A4E1D15035B283D3FDF616CC (I2F2159E4520CF0D6E57382C8E60EC46D ),
.I2EF8304B3AEA32E6C6F568223FAD9CBA (IC1C88613A52A238F417438A678D1196A ), .I369C6CA451B73B45E1F8D4D8AA53C2AD (I673AF3DF8D93FAFCF8E255C8C6852D9B ),
.IE81278F89BAA90C1F6EF0784D0DE2F62 (I2BE5B3BCC47A675D856661ED2CA18C19 ), .I2F86B5F8620848A51ED4F1F736CF8825 (I4DDF7CB99428D62C1FB17E5C8FA42E6A ),
.I63FDDFAA5AB093F3BB343A8C133F3BAF (I7B40A3A5ECAB9C16D0C5E2614F94A037 ), .IE7F8A35B24BC8805CAD86FD378C18296 (IB76DC52DFFF4905395FBC5C33F2C6B24 ),
.IAB90D3559ED5004EBCCD9D73A2928E3F (I8236407E542CBF20A06054E415DF3019 ), .I75EB9BE30F2D20C56659251E3B505209 (I45B614E1199C70B4E5F58D3EFD1D08C7 ),
.I3E8F0524CDEE96F573376A6BF670184B (I69B84382CF4434D3BBB964B953CD6E15 ), .I17066520A25539E7F98555DFF7832BBE (IF66089F4B958743DD8052C5F9D832CD1 ),
.IB33B8D629A269D1BC3D79902EE2EB312 (IA69B6A69D96E898639A555BF6567C273 ), .I1E494BBA2ECB063404DBB73667CC7E8D (IFD8A5AA76F99D6914AE0274FCD000AD1 ),
.I4A4976CAF016EA789DCDB7AA131246C3 (ICA6FC4E4455EED217775291436AD860C ), .I5ADFC7E7F8B570F5258C2813D0020950 (IFE46A9371C863D1229E8DCA840188E17 ),
.I1FD27F5D298FA5493F3F510610F19E4E (IF63E39473014C2B5C4FB8832104F3754 ), .IEA9D116BFADD4042E3D3AD0C618B652A (I58FB5703785F6B602E564F2C3886577D ),
.I418D7ADEC09B065FFE6565D649D285B6 (IC85FD97ECAC87466B9C19ACECC79FC2D ), .IF2B42773D268BA706D29FCCFCB799AF9 (IA5B538B804B78BFE2529013B5C97D493 ),
.I470C1C74A2768E559679EE12280C8506 (IB7543BE04BDCE5E5193E442BACB25B09 ), .I513461A4DA46CAA79BEC76A8DE8E2A98 (IC6D81493F78B34E8262D34CE51650B27 ),
.ID7F4713F32DABD57E54222A946FA802F (ID40108F42D0FA32BFA839EFAD8F8C320 ), .IADE62F3832E7DA9091E0F5B2EBC50F9C (I46618BF7FF1CE70399E81FFAD2D6846B ),
.I3443654006276E8DC7EE67AAE2283C64 (I1CA27197DF7539251654AB3DAC8E8B38 ), .I4FD27244D7DB92B0548A7AE35BDEDE28 (I755156D55303F238FD088C21A8C23864 ),
.IDB44E9A441DC017FFA044AB8E232791F (ID2C4F123A6A9197C7B4B4FD780FCC272 ) ); end endgenerate ICF327C89C36124513E146F1FF3BCDEEB
#( .I87C69AEB153025D890F0A7CE399F00FE (IBACE8243A55E1A6C355E86BA25034EFB ), .I68B4790A0165FFB6E2740B409126FE6B (8),
.I66C185998F46A7148163982E39BCD296 (I66C185998F46A7148163982E39BCD296 ) )  IA440041682C400211AAD0D987978451E ( .ICCFB0F435B37370076102F325BC08D20
(ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .I0C5BEBB297319D36CFD96B791AFE888C
(ID2C4F123A6A9197C7B4B4FD780FCC272 ), .I42D2723FE4CDE4AF565DD01BD32BB8AC (I42D2723FE4CDE4AF565DD01BD32BB8AC ), .I8E99DEF5C63C6A55606BD30E4BE8E3FB
(I8E99DEF5C63C6A55606BD30E4BE8E3FB ), .IC3760F6E74F9AA61561390CC1466FC1A (IC3760F6E74F9AA61561390CC1466FC1A ), .I582940C94DBA710A62923187D833E8E6
(I582940C94DBA710A62923187D833E8E6 ), .IAFF3235BDF22DE6B7D7DBF12451FA2FE (I48ABEC51DF27ACA5596235F4DF0D08C4 ), .I5FFD1878342C11E50C1617928EBB38D7
(IF77AAC35DEF2E12949B516C97BABF4FD ), .I27766E6DFBDE7E37CDB16F4E2C0E1DD4 (I586E9AE745283DB69A128B0C7A472DE0 ), .I520751EAD225B5BFC3D7E0ACB7BC6405
(I91383F42CED2732A542098CD5ACFFD1D ), .IFA5857E29877E868702F9890224BA5FC (I45B614E1199C70B4E5F58D3EFD1D08C7 ), .I3CEE775C269D38D2B516507E40A6387C
(I69B84382CF4434D3BBB964B953CD6E15 ), .IEADE52DA6BAC6B55AC606944635D8C9A (IF66089F4B958743DD8052C5F9D832CD1 ) );
I6433000F3EF06E04177C32D16C534889 # ( .IB71844FFA3AB85FEF45EAB4D35395752 (I99651B9F47529E0ADC5349B57C84E531 ), .I5C6C6CD7723900C21B3A76E887CEE164
(I6684631E4DAAC3FB7551EF267A7E3D73 ), .I64BB723AC8F87F7AEBA73BF190ED5F8F (I7292F55C07BFD7FB8A60D29FFC186275 ), .I66C185998F46A7148163982E39BCD296
(I66C185998F46A7148163982E39BCD296 ) )  I4FE5E72F36162FB85A7454C2F371EED7 ( .ICCFB0F435B37370076102F325BC08D20 (ICCFB0F435B37370076102F325BC08D20 ),
.I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .I27CF4DD7FCBC7E0A229344EDF94F2651 (I58FB5703785F6B602E564F2C3886577D ),
.I1A55EB74BDB9184AA980B07905C85479 (IC85FD97ECAC87466B9C19ACECC79FC2D ), .I48D61F5A0B5732A58912433B42CD9D0C (ID40108F42D0FA32BFA839EFAD8F8C320 ),
.I04BC24D2B6403E54A64DE9E6C9ABAA2B (I884F4ADE09FABBA20600F67BC1A50FE7 ), .I3F6FB755DC9826D564C143FF9E32F032 (I61E8E6981294A3342BDF5596043A2DFA ),
.IE315CDCA06C9620D5C0AB966E553F0C3 (I2F5C52C0CABA5EFAF34A96BC39DA8F96 ), .ID7FCE45A65ADDB17F91F73A1B506BB5B ( ),
.I125028C7446331521D0434C10E8B0007 (I2F2159E4520CF0D6E57382C8E60EC46D ), .I8BB939FF2AFDE7B2A1E480DCB61CE354 (I4DDF7CB99428D62C1FB17E5C8FA42E6A ),
.IC9DE8233C6B1ADF4418EEF5B1F14BE49 (IA4EA76535E7026B1F7DF3EDC236AF756 ), .I585F74DE05DD9C1C7070D6B4F6E181C2 (I7DA036F5B0B44A1D5E3EB0237828A810 ),
.I233E0C0C8E5150F0CD8258F276D93942 (I7F72A1B5D33702E3B645BD20CB425937 ), .IBE0D6810EBD63B5C428623C578CF6D3A ( )
); I6433000F3EF06E04177C32D16C534889 # ( .IB71844FFA3AB85FEF45EAB4D35395752 (I0AEF008AE3BC7E23C49F86BC2B344750 ),
.I5C6C6CD7723900C21B3A76E887CEE164 (I6684631E4DAAC3FB7551EF267A7E3D73 ), .I64BB723AC8F87F7AEBA73BF190ED5F8F (I7292F55C07BFD7FB8A60D29FFC186275 ),
.I66C185998F46A7148163982E39BCD296 (I66C185998F46A7148163982E39BCD296 ) )  I48BFA8FF344ECC3BA7AAD048A7985C79 ( .ICCFB0F435B37370076102F325BC08D20
(ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .I27CF4DD7FCBC7E0A229344EDF94F2651
(I58FB5703785F6B602E564F2C3886577D ), .I1A55EB74BDB9184AA980B07905C85479 (IB7543BE04BDCE5E5193E442BACB25B09 ), .I48D61F5A0B5732A58912433B42CD9D0C
(I1CA27197DF7539251654AB3DAC8E8B38 ), .I04BC24D2B6403E54A64DE9E6C9ABAA2B (IA5896E672427191F9A0B4ED1C9301313 ), .I3F6FB755DC9826D564C143FF9E32F032
(I0317313DEECD8AC19E98BA2F1C27E0A9 ), .IE315CDCA06C9620D5C0AB966E553F0C3 (IFDB2ACAC637F40CDDFBB20A3AFD9A401 ), .ID7FCE45A65ADDB17F91F73A1B506BB5B
( ), .I125028C7446331521D0434C10E8B0007 (I673AF3DF8D93FAFCF8E255C8C6852D9B ), .I8BB939FF2AFDE7B2A1E480DCB61CE354
(IB76DC52DFFF4905395FBC5C33F2C6B24 ), .IC9DE8233C6B1ADF4418EEF5B1F14BE49 (I9D0CEC2083A8932FA283AD091303049F ), .I585F74DE05DD9C1C7070D6B4F6E181C2
(IE43DA634E45C0D88369455568042AF37 ), .I233E0C0C8E5150F0CD8258F276D93942 (IB6FE1681C40869E515EA3BF2BD5F7DA8 ), .IBE0D6810EBD63B5C428623C578CF6D3A
( ) ); I6433000F3EF06E04177C32D16C534889 # ( .IB71844FFA3AB85FEF45EAB4D35395752 (I0AEF008AE3BC7E23C49F86BC2B344750 ),
.I5C6C6CD7723900C21B3A76E887CEE164 (I3A59A966031A54015DBF77A68A5A82D3 ), .I64BB723AC8F87F7AEBA73BF190ED5F8F (I7292F55C07BFD7FB8A60D29FFC186275 ),
.I66C185998F46A7148163982E39BCD296 (I66C185998F46A7148163982E39BCD296 ) )  IC6BE0D645D48779DADE25A4973891991 ( .ICCFB0F435B37370076102F325BC08D20
(ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .I27CF4DD7FCBC7E0A229344EDF94F2651
(I58FB5703785F6B602E564F2C3886577D ), .I1A55EB74BDB9184AA980B07905C85479 (IC6D81493F78B34E8262D34CE51650B27 ), .I48D61F5A0B5732A58912433B42CD9D0C
(I755156D55303F238FD088C21A8C23864 ), .I04BC24D2B6403E54A64DE9E6C9ABAA2B (IE4C3654339F6BF285840C2AB868371A1 ), .I3F6FB755DC9826D564C143FF9E32F032
(I5F40D6DD3270B21E2E90925F127E6477 ), .IE315CDCA06C9620D5C0AB966E553F0C3 (I33A8C146E90D24E54E605500849CD461 ), .ID7FCE45A65ADDB17F91F73A1B506BB5B
( ), .I125028C7446331521D0434C10E8B0007 (I2BE5B3BCC47A675D856661ED2CA18C19 ), .I8BB939FF2AFDE7B2A1E480DCB61CE354
(I8236407E542CBF20A06054E415DF3019 ), .IC9DE8233C6B1ADF4418EEF5B1F14BE49 (I173FA018899178893FB946275729ED68 ), .I585F74DE05DD9C1C7070D6B4F6E181C2
(I5871F7D82773EB9D3EE955FCC1611D9F ), .I233E0C0C8E5150F0CD8258F276D93942 (I96EC08C26A305FC6029163D693EF44E6 ), .IBE0D6810EBD63B5C428623C578CF6D3A
( ) ); I6433000F3EF06E04177C32D16C534889 # ( .IB71844FFA3AB85FEF45EAB4D35395752 (ICED1C5B792370B25488CFA18FE5E472E ),
.I5C6C6CD7723900C21B3A76E887CEE164 (I3A59A966031A54015DBF77A68A5A82D3 ), .I64BB723AC8F87F7AEBA73BF190ED5F8F (I7292F55C07BFD7FB8A60D29FFC186275 ),
.I66C185998F46A7148163982E39BCD296 (I66C185998F46A7148163982E39BCD296 ) )  IDFB6DB2CA10C61E108DCCB4FB9528FEB ( .ICCFB0F435B37370076102F325BC08D20
(ICCFB0F435B37370076102F325BC08D20 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7 (I9ED2A9117D3AEAF54CBA7AD69083BCB7 ), .I27CF4DD7FCBC7E0A229344EDF94F2651
(I58FB5703785F6B602E564F2C3886577D ), .I1A55EB74BDB9184AA980B07905C85479 (IA5B538B804B78BFE2529013B5C97D493 ), .I48D61F5A0B5732A58912433B42CD9D0C
(I46618BF7FF1CE70399E81FFAD2D6846B ), .I04BC24D2B6403E54A64DE9E6C9ABAA2B (I0BA940AC86B853EFCE63667C128E2DF4 ), .I3F6FB755DC9826D564C143FF9E32F032
(ID176017A6F96653AFD707B70D22BEA8C ), .IE315CDCA06C9620D5C0AB966E553F0C3 (IE8C34BE7792A66A23CB1C7A5CFF55BBF ), .ID7FCE45A65ADDB17F91F73A1B506BB5B
( ), .I125028C7446331521D0434C10E8B0007 (IC1C88613A52A238F417438A678D1196A ), .I8BB939FF2AFDE7B2A1E480DCB61CE354
(I7B40A3A5ECAB9C16D0C5E2614F94A037 ), .IC9DE8233C6B1ADF4418EEF5B1F14BE49 (ID505752183B05B70B86F1045E7DB0CF0 ), .I585F74DE05DD9C1C7070D6B4F6E181C2
(I36AD11753E1A0E22546912955186E616 ), .I233E0C0C8E5150F0CD8258F276D93942 (I5E12F1044C6612C74B661A7400A97D4B ), .IBE0D6810EBD63B5C428623C578CF6D3A
( ) ); endmodule 
  module pcie_mfdev_subsys #( parameter gx_cs_f0_bar0_size = "NONE", gx_cs_f0_bar0_is_64_bit = 0, gx_cs_f0_bar0_is_io_space
= 0, gx_cs_f0_bar0_is_prefetchable = 1, gx_cs_f0_bar1_size = "NONE", gx_cs_f0_bar1_is_io_space = 0, gx_cs_f0_bar1_is_prefetchable
= 1, gx_cs_f0_bar2_size = "NONE", gx_cs_f0_bar2_is_64_bit = 0, gx_cs_f0_bar2_is_io_space = 0, gx_cs_f0_bar2_is_prefetchable
= 1, gx_cs_f0_bar3_size = "NONE", gx_cs_f0_bar3_is_io_space = 0, gx_cs_f0_bar3_is_prefetchable = 1, gx_cs_f0_bar4_size
= "NONE", gx_cs_f0_bar4_is_64_bit = 0, gx_cs_f0_bar4_is_io_space = 0, gx_cs_f0_bar4_is_prefetchable = 1, gx_cs_f0_bar5_size
= "NONE", gx_cs_f0_bar5_is_io_space = 0, gx_cs_f0_bar5_is_prefetchable = 1, gx_cs_f0_class_code = 24'h000000, gx_cs_f0_device_id
= 16'h0000, gx_cs_f0_int_count = 1, gx_cs_f0_int_pin = "INTA", gx_cs_f0_revision_id = 8'h00, gx_cs_f0_subsystem_id
= 16'h0000, gx_cs_f1_bar0_size = "NONE", gx_cs_f1_bar0_is_64_bit = 0, gx_cs_f1_bar0_is_io_space = 0, gx_cs_f1_bar0_is_prefetchable
= 1, gx_cs_f1_bar1_size = "NONE", gx_cs_f1_bar1_is_io_space = 0, gx_cs_f1_bar1_is_prefetchable = 1, gx_cs_f1_bar2_size
= "NONE", gx_cs_f1_bar2_is_64_bit = 0, gx_cs_f1_bar2_is_io_space = 0, gx_cs_f1_bar2_is_prefetchable = 1, gx_cs_f1_bar3_size
= "NONE", gx_cs_f1_bar3_is_io_space = 0, gx_cs_f1_bar3_is_prefetchable = 1, gx_cs_f1_bar4_size = "NONE", gx_cs_f1_bar4_is_64_bit
= 0, gx_cs_f1_bar4_is_io_space = 0, gx_cs_f1_bar4_is_prefetchable = 1, gx_cs_f1_bar5_size = "NONE", gx_cs_f1_bar5_is_io_space
= 0, gx_cs_f1_bar5_is_prefetchable = 1, gx_cs_f1_class_code = 24'h000000, gx_cs_f1_device_id = 16'h0000, gx_cs_f1_int_count
= 0, gx_cs_f1_int_pin = "INTA", gx_cs_f1_present = 0, gx_cs_f1_revision_id = 8'h00, gx_cs_f1_subsystem_id = 16'h0000,
gx_cs_f2_bar0_size = "NONE", gx_cs_f2_bar0_is_64_bit = 0, gx_cs_f2_bar0_is_io_space = 0, gx_cs_f2_bar0_is_prefetchable
= 1, gx_cs_f2_bar1_size = "NONE", gx_cs_f2_bar1_is_io_space = 0, gx_cs_f2_bar1_is_prefetchable = 1, gx_cs_f2_bar2_size
= "NONE", gx_cs_f2_bar2_is_64_bit = 0, gx_cs_f2_bar2_is_io_space = 0, gx_cs_f2_bar2_is_prefetchable = 1, gx_cs_f2_bar3_size
= "NONE", gx_cs_f2_bar3_is_io_space = 0, gx_cs_f2_bar3_is_prefetchable = 1, gx_cs_f2_bar4_size = "NONE", gx_cs_f2_bar4_is_64_bit
= 0, gx_cs_f2_bar4_is_io_space = 0, gx_cs_f2_bar4_is_prefetchable = 1, gx_cs_f2_bar5_size = "NONE", gx_cs_f2_bar5_is_io_space
= 0, gx_cs_f2_bar5_is_prefetchable = 1, gx_cs_f2_class_code = 24'h000000, gx_cs_f2_device_id = 16'h0000, gx_cs_f2_int_count
= 0, gx_cs_f2_int_pin = "INTA", gx_cs_f2_present = 0, gx_cs_f2_revision_id = 8'h00, gx_cs_f2_subsystem_id = 16'h0000,
gx_cs_f3_bar0_size = "NONE", gx_cs_f3_bar0_is_64_bit = 0, gx_cs_f3_bar0_is_io_space = 0, gx_cs_f3_bar0_is_prefetchable
= 1, gx_cs_f3_bar1_size = "NONE", gx_cs_f3_bar1_is_io_space = 0, gx_cs_f3_bar1_is_prefetchable = 1, gx_cs_f3_bar2_size
= "NONE", gx_cs_f3_bar2_is_64_bit = 0, gx_cs_f3_bar2_is_io_space = 0, gx_cs_f3_bar2_is_prefetchable = 1, gx_cs_f3_bar3_size
= "NONE", gx_cs_f3_bar3_is_io_space = 0, gx_cs_f3_bar3_is_prefetchable = 1, gx_cs_f3_bar4_size = "NONE", gx_cs_f3_bar4_is_64_bit
= 0, gx_cs_f3_bar4_is_io_space = 0, gx_cs_f3_bar4_is_prefetchable = 1, gx_cs_f3_bar5_size = "NONE", gx_cs_f3_bar5_is_io_space
= 0, gx_cs_f3_bar5_is_prefetchable = 1, gx_cs_f3_class_code = 24'h000000, gx_cs_f3_device_id = 16'h0000, gx_cs_f3_int_count
= 0, gx_cs_f3_int_pin = "INTA", gx_cs_f3_present = 0, gx_cs_f3_revision_id = 8'h00, gx_cs_f3_subsystem_id = 16'h0000,
gx_cs_f4_bar0_size = "NONE", gx_cs_f4_bar0_is_64_bit = 0, gx_cs_f4_bar0_is_io_space = 0, gx_cs_f4_bar0_is_prefetchable
= 1, gx_cs_f4_bar1_size = "NONE", gx_cs_f4_bar1_is_io_space = 0, gx_cs_f4_bar1_is_prefetchable = 1, gx_cs_f4_bar2_size
= "NONE", gx_cs_f4_bar2_is_64_bit = 0, gx_cs_f4_bar2_is_io_space = 0, gx_cs_f4_bar2_is_prefetchable = 1, gx_cs_f4_bar3_size
= "NONE", gx_cs_f4_bar3_is_io_space = 0, gx_cs_f4_bar3_is_prefetchable = 1, gx_cs_f4_bar4_size = "NONE", gx_cs_f4_bar4_is_64_bit
= 0, gx_cs_f4_bar4_is_io_space = 0, gx_cs_f4_bar4_is_prefetchable = 1, gx_cs_f4_bar5_size = "NONE", gx_cs_f4_bar5_is_io_space
= 0, gx_cs_f4_bar5_is_prefetchable = 1, gx_cs_f4_class_code = 24'h000000, gx_cs_f4_device_id = 16'h0000, gx_cs_f4_int_count
= 0, gx_cs_f4_int_pin = "INTA", gx_cs_f4_present = 0, gx_cs_f4_revision_id = 8'h00, gx_cs_f4_subsystem_id = 16'h0000,
gx_cs_f5_bar0_size = "NONE", gx_cs_f5_bar0_is_64_bit = 0, gx_cs_f5_bar0_is_io_space = 0, gx_cs_f5_bar0_is_prefetchable
= 1, gx_cs_f5_bar1_size = "NONE", gx_cs_f5_bar1_is_io_space = 0, gx_cs_f5_bar1_is_prefetchable = 1, gx_cs_f5_bar2_size
= "NONE", gx_cs_f5_bar2_is_64_bit = 0, gx_cs_f5_bar2_is_io_space = 0, gx_cs_f5_bar2_is_prefetchable = 1, gx_cs_f5_bar3_size
= "NONE", gx_cs_f5_bar3_is_io_space = 0, gx_cs_f5_bar3_is_prefetchable = 1, gx_cs_f5_bar4_size = "NONE", gx_cs_f5_bar4_is_64_bit
= 0, gx_cs_f5_bar4_is_io_space = 0, gx_cs_f5_bar4_is_prefetchable = 1, gx_cs_f5_bar5_size = "NONE", gx_cs_f5_bar5_is_io_space
= 0, gx_cs_f5_bar5_is_prefetchable = 1, gx_cs_f5_class_code = 24'h000000, gx_cs_f5_device_id = 16'h0000, gx_cs_f5_int_count
= 0, gx_cs_f5_int_pin = "INTA", gx_cs_f5_present = 0, gx_cs_f5_revision_id = 8'h00, gx_cs_f5_subsystem_id = 16'h0000,
gx_cs_f6_bar0_size = "NONE", gx_cs_f6_bar0_is_64_bit = 0, gx_cs_f6_bar0_is_io_space = 0, gx_cs_f6_bar0_is_prefetchable
= 1, gx_cs_f6_bar1_size = "NONE", gx_cs_f6_bar1_is_io_space = 0, gx_cs_f6_bar1_is_prefetchable = 1, gx_cs_f6_bar2_size
= "NONE", gx_cs_f6_bar2_is_64_bit = 0, gx_cs_f6_bar2_is_io_space = 0, gx_cs_f6_bar2_is_prefetchable = 1, gx_cs_f6_bar3_size
= "NONE", gx_cs_f6_bar3_is_io_space = 0, gx_cs_f6_bar3_is_prefetchable = 1, gx_cs_f6_bar4_size = "NONE", gx_cs_f6_bar4_is_64_bit
= 0, gx_cs_f6_bar4_is_io_space = 0, gx_cs_f6_bar4_is_prefetchable = 1, gx_cs_f6_bar5_size = "NONE", gx_cs_f6_bar5_is_io_space
= 0, gx_cs_f6_bar5_is_prefetchable = 1, gx_cs_f6_class_code = 24'h000000, gx_cs_f6_device_id = 16'h0000, gx_cs_f6_int_count
= 0, gx_cs_f6_int_pin = "INTA", gx_cs_f6_present = 0, gx_cs_f6_revision_id = 8'h00, gx_cs_f6_subsystem_id = 16'h0000,
gx_cs_f7_bar0_size = "NONE", gx_cs_f7_bar0_is_64_bit = 0, gx_cs_f7_bar0_is_io_space = 0, gx_cs_f7_bar0_is_prefetchable
= 1, gx_cs_f7_bar1_size = "NONE", gx_cs_f7_bar1_is_io_space = 0, gx_cs_f7_bar1_is_prefetchable = 1, gx_cs_f7_bar2_size
= "NONE", gx_cs_f7_bar2_is_64_bit = 0, gx_cs_f7_bar2_is_io_space = 0, gx_cs_f7_bar2_is_prefetchable = 1, gx_cs_f7_bar3_size
= "NONE", gx_cs_f7_bar3_is_io_space = 0, gx_cs_f7_bar3_is_prefetchable = 1, gx_cs_f7_bar4_size = "NONE", gx_cs_f7_bar4_is_64_bit
= 0, gx_cs_f7_bar4_is_io_space = 0, gx_cs_f7_bar4_is_prefetchable = 1, gx_cs_f7_bar5_size = "NONE", gx_cs_f7_bar5_is_io_space
= 0, gx_cs_f7_bar5_is_prefetchable = 1, gx_cs_f7_class_code = 24'h000000, gx_cs_f7_device_id = 16'h0000, gx_cs_f7_int_count
= 0, gx_cs_f7_int_pin = "INTA", gx_cs_f7_present = 0, gx_cs_f7_revision_id = 8'h00, gx_cs_f7_subsystem_id = 16'h0000,
gx_cs_subsystem_vendor_id = 16'h0000, gx_cs_vendor_id = 16'h0000, gx_ipx_data_sz = 16, gx_nr_wb_tgts = 3, gx_pcie_gen2
= 0, gx_tech_lib = "ECP3", gx_wbm_data_sz = 32, gx_wbs_data_sz = 32, gx_wbm_adr_sz = 24, gx_wbs_adr_sz = 48 ) (
input wire ix_clk_125 ,  input wire ix_rst_n , input wire [gx_nr_wb_tgts - 1:0] ix_dec_wb_cyc , input wire ix_ipx_dl_up ,
input wire ix_ipx_malf_tlp , input wire [2:0] ix_ipx_pcie_linkw , input wire ix_ipx_pcie_rate , input wire [gx_ipx_data_sz
- 1:0] ix_ipx_rx_data , input wire ix_ipx_rx_dwen , input wire ix_ipx_rx_end , input wire ix_ipx_rx_st , input wire
[12:0] ix_ipx_tx_ca_cpld , input wire [8:0] ix_ipx_tx_ca_cplh , input wire [12:0] ix_ipx_tx_ca_npd , input wire
[8:0] ix_ipx_tx_ca_nph , input wire [12:0] ix_ipx_tx_ca_pd , input wire [8:0] ix_ipx_tx_ca_ph , input wire ix_ipx_tx_rdy ,
input wire ix_ipx_tx_val , input wire [gx_cs_f7_int_count + gx_cs_f6_int_count + gx_cs_f5_int_count + gx_cs_f4_int_count
+ gx_cs_f3_int_count + gx_cs_f2_int_count + gx_cs_f1_int_count + gx_cs_f0_int_count - 1:0] ix_pci_int_req , input
wire [31:0] ix_pci_rsz_f0_bar0 ,  input wire [31:0] ix_pci_rsz_f0_bar1 , input wire [31:0] ix_pci_rsz_f0_bar2 ,
input wire [31:0] ix_pci_rsz_f0_bar3 , input wire [31:0] ix_pci_rsz_f0_bar4 , input wire [31:0] ix_pci_rsz_f0_bar5 ,
input wire [31:0] ix_pci_rsz_f1_bar0 , input wire [31:0] ix_pci_rsz_f1_bar1 , input wire [31:0] ix_pci_rsz_f1_bar2 ,
input wire [31:0] ix_pci_rsz_f1_bar3 , input wire [31:0] ix_pci_rsz_f1_bar4 , input wire [31:0] ix_pci_rsz_f1_bar5 ,
input wire [31:0] ix_pci_rsz_f2_bar0 , input wire [31:0] ix_pci_rsz_f2_bar1 , input wire [31:0] ix_pci_rsz_f2_bar2 ,
input wire [31:0] ix_pci_rsz_f2_bar3 , input wire [31:0] ix_pci_rsz_f2_bar4 , input wire [31:0] ix_pci_rsz_f2_bar5 ,
input wire [31:0] ix_pci_rsz_f3_bar0 , input wire [31:0] ix_pci_rsz_f3_bar1 , input wire [31:0] ix_pci_rsz_f3_bar2 ,
input wire [31:0] ix_pci_rsz_f3_bar3 , input wire [31:0] ix_pci_rsz_f3_bar4 , input wire [31:0] ix_pci_rsz_f3_bar5 ,
input wire [31:0] ix_pci_rsz_f4_bar0 , input wire [31:0] ix_pci_rsz_f4_bar1 , input wire [31:0] ix_pci_rsz_f4_bar2 ,
input wire [31:0] ix_pci_rsz_f4_bar3 , input wire [31:0] ix_pci_rsz_f4_bar4 , input wire [31:0] ix_pci_rsz_f4_bar5 ,
input wire [31:0] ix_pci_rsz_f5_bar0 , input wire [31:0] ix_pci_rsz_f5_bar1 , input wire [31:0] ix_pci_rsz_f5_bar2 ,
input wire [31:0] ix_pci_rsz_f5_bar3 , input wire [31:0] ix_pci_rsz_f5_bar4 , input wire [31:0] ix_pci_rsz_f5_bar5 ,
input wire [31:0] ix_pci_rsz_f6_bar0 , input wire [31:0] ix_pci_rsz_f6_bar1 , input wire [31:0] ix_pci_rsz_f6_bar2 ,
input wire [31:0] ix_pci_rsz_f6_bar3 , input wire [31:0] ix_pci_rsz_f6_bar4 , input wire [31:0] ix_pci_rsz_f6_bar5 ,
input wire [31:0] ix_pci_rsz_f7_bar0 , input wire [31:0] ix_pci_rsz_f7_bar1 , input wire [31:0] ix_pci_rsz_f7_bar2 ,
input wire [31:0] ix_pci_rsz_f7_bar3 , input wire [31:0] ix_pci_rsz_f7_bar4 , input wire [31:0] ix_pci_rsz_f7_bar5 ,
input wire ix_wbm_ack , input wire [gx_wbm_data_sz - 1:0] ix_wbm_dat , input wire ix_wbm_err , input wire [gx_wbs_adr_sz
- 1:0] ix_wbs_adr , input wire [1:0] ix_wbs_bte , input wire [2:0] ix_wbs_cti , input wire [7:0] ix_wbs_cyc , input
wire [gx_wbs_data_sz - 1:0] ix_wbs_dat , input wire [(gx_wbs_data_sz / 8) - 1:0] ix_wbs_sel , input wire ix_wbs_stb ,
input wire ix_wbs_we , output wire [gx_wbm_adr_sz - 1:0] ox_dec_adr , output wire [5:0] ox_dec_bar_hit , output
wire [7:0] ox_dec_func_hit , output wire [7:0] ox_ipx_cc_npd_num , output wire [7:0] ox_ipx_cc_pd_num , output wire
ox_ipx_cc_processed_npd , output wire ox_ipx_cc_processed_nph , output wire ox_ipx_cc_processed_pd , output wire
ox_ipx_cc_processed_ph , output wire [gx_ipx_data_sz - 1:0] ox_ipx_tx_data , output wire ox_ipx_tx_dwen , output
wire ox_ipx_tx_end , output wire ox_ipx_tx_req , output wire ox_ipx_tx_st , output wire [gx_wbm_adr_sz - 1:0] ox_wbm_adr ,
output wire [1:0] ox_wbm_bte , output wire [2:0] ox_wbm_cti , output wire [gx_nr_wb_tgts - 1:0] ox_wbm_cyc , output
wire [gx_wbm_data_sz - 1:0] ox_wbm_dat , output wire [(gx_wbm_data_sz / 8) - 1:0] ox_wbm_sel , output wire ox_wbm_stb ,
output wire ox_wbm_we , output wire ox_wbs_ack , output wire [gx_wbs_data_sz - 1:0] ox_wbs_dat , output wire ox_wbs_err ,
output wire ox_sys_rst_n , output wire [7:0] ox_sys_rst_func_n );   localparam IEF532EA44160288B0ED6812C670E4CDB
= gx_wbm_data_sz ; localparam I96690071F3CE4794E376870D1BB87C22 = (gx_ipx_data_sz == 16) ? 32 : 64; localparam I249BB13F12A1B213E14013F118AB1013
= I96690071F3CE4794E376870D1BB87C22 / gx_wbm_data_sz ; localparam I37BDD1A019498B0050A3FF971DCE0165 = (gx_ipx_data_sz
> gx_wbm_data_sz ) ? 1 : 0; localparam I90D984439DDA58639C67AC709C0E6CC9 = 1024;  localparam IC6E51C590A86FEEF8592133ED3A689E7
= $clog2((I90D984439DDA58639C67AC709C0E6CC9 * I249BB13F12A1B213E14013F118AB1013 ) + 1); localparam I31F00D08C3CE05C5A25E18130CAFEAD5
= 512;  localparam I9A19F862D1FD27BAC93F9AC85F8F1B2B = $clog2((I31F00D08C3CE05C5A25E18130CAFEAD5 * I249BB13F12A1B213E14013F118AB1013 )
+ 1); localparam I51E5032D35684B1A6595F2291E95EBFD = 512;  localparam IB985C42C0963EF96E8DAFEE1BF657C01 = $clog2((I51E5032D35684B1A6595F2291E95EBFD
* I249BB13F12A1B213E14013F118AB1013 ) + 1); localparam IF3D376C350B88011F1FC2F939263D178 = 512;  localparam I8224701A907960C6458368B9E178E270
= $clog2((IF3D376C350B88011F1FC2F939263D178 * I249BB13F12A1B213E14013F118AB1013 ) + 1); localparam IB89F6B40906A7C6F23E0C9CD1176DAD6
= 1024;  localparam I7C43BE354681C8AAA7229179D47CE564 = $clog2(IB89F6B40906A7C6F23E0C9CD1176DAD6 + 1); localparam
IB18B8E96B09D7E54E97338C01ECBF348 = (gx_wbm_adr_sz < 15) ? 15 : gx_wbm_adr_sz ;  wire IB552918C70C5F8374FC906E0C2225F89 ;
wire [I96690071F3CE4794E376870D1BB87C22 - 1:0] IE593D61A89622FBF1D4D61DBF77B0759 ; wire IEB0657AD1CF8431866F1DACFA91DAE9C ;
wire I09D474E43198BB26D683E473E35C90C8 ; wire IA51154D40B341A92D3FF48956FE47EDD ; wire [I7C43BE354681C8AAA7229179D47CE564
- 1:0] I2FB68C8CAC3EE2BC47F461C034FBC722 ; wire [IEF532EA44160288B0ED6812C670E4CDB - 1:0] I78FE781BC8B5C49E9E0559250B6D4289 ;
wire IA5B0FE243F631FAA054C108CC3F72E10 ; wire IE228EF2D803387145092976501986E10 ; wire I6DF8AFD2D5E8EFB85D4507AC54B8E25C ;
wire [7:0] IF60FDFFF213C716383F950A9422A1758 ; wire [7:0] I4FF065235743696A883B835CA5B1B85D ; wire IA4F8AA6824642C6A9DC9A7747287580D ;
wire I010A8CBEA176E0F2178CBA8B77E6FE07 ; wire I00B00319AA148C3D5F9C641ABDDBAFA3 ; wire I92625F81A8AD6C4657526FD7E7F0D00C ;
wire [63:0] I220A96CF74656D5120C8D113E4B1ED55 ; wire IBE8D7D536CBDF087E7E00B93DA215E3D ; wire I4DC446D96F0774A667A70D52D9392874 ;
wire I3FF9BAFBF91288E78D7EA6DD95DB3A40 ; wire [7:0] IE67E5659AC07E2D371890CDACFA6ED42 ; wire [4:0] I18137FEBF7FA4CE04FDE793386121F57 ;
wire [2:0] I0B37325C0AB5EEA3148286371EB202D1 ; wire IAF786EDCB7BC54665688D1FC2E0E922F ; wire [IEF532EA44160288B0ED6812C670E4CDB
- 1:0] I6609F40DB9BF2AAD262974646AD5EBE5 ; wire IAE96F702FDFFAF4D7DD2303A7E5CAA82 ; wire I314F20E260B367A911975FFD9E094426 ;
wire I4A399AD6EACAD372F1F0ED553AF29E10 ; wire [IB18B8E96B09D7E54E97338C01ECBF348 - 1:0] IE81C89DB2F6C737F2D82BE35AFC7DDA2 ;
wire [1:0] IC13572948B0A4216A965E35100DE669F ; wire [2:0] I599F86FA1B9AEED5B32EE8B27DFFFACE ; wire I291FF0AF6B998FB4D8BD958CFDA1CF8C ;
wire [gx_nr_wb_tgts - 1: 0] IDCB78AD56EF8FEF35AAF4DED8D1F87B6 ; wire [gx_wbm_data_sz - 1:0] IEC017B3AB9F16AE871D5253A5257D941 ;
wire [3:0] I87343FD56CEFDCB10F9A272CF1F0CA8E ; wire IB8F3718FAD7719FD71FDE3B0DE8D7445 ; wire IB6F57A3FE1F5B6A182168AC92AC3D457 ;
wire [10:0] I7681E0E609A03559F13166ACF7852905 ; wire [3:0] I507A0A1A3C69E79845F5C15AFFAF6595 ; wire [3:0] IDB0B420EA96A60B402FECD3AE3620DCC ;
wire I678B3227DE7FFEFE726CE68123B91F8D ; wire [7:0] I4BA2D171F5FD7E0FEACB9DF4C87DDC19 ; wire IC0197882115D001485B37646159E234E ;
wire [7:0] IB1AAAED8469CADFA3AB4BF806A8466B6 ; wire IA6774F4F4F3AF83C6A9E233DB00F89A0 ; wire IFFF50035216FD68A74F8164F0EE74689 ;
wire IF9A16909C25386742335A246DEDE12E8 ; wire I5078F81AE0F5DCD4CC2ABEE2CEF9C827 ; wire IB55475954FE95F83F22B1C2FB76FAEC7 ;
wire I31980ABC07D19BA89784085C7754DE42 ; wire [7:0] IE1F9397E899B4E938A0D54FC51445C13 ; wire [2:0] IDE0F2D42601304C0E0CCD60778B3938F ;
wire [7:0] I395C5996AD91572D0F6652373B6018E7 ; wire [4:0] I5B507E107F91FDBF0B2EEF7DD9AE40C5 ; wire [2:0] IBAE868C7DE15BF2F751B0177B798BDCD ;
wire [2:0] IAF2A92B584FD036A9F751EB8F3FA7ACD ; wire [2:0] I5CF35907FA895D81AAC1AAFED86DBE1F ; wire [7:0] I1BAAE01807D45E9F21D2ACB2BCB4F621 ;
wire ID872B1CCC580E5915A782E136C7A691B ; wire [31:0] IFFB9EED620356BDFB94697DB3606174F ; wire I2C072E656BFCADF4877B42244D6D2307 ;
wire IB96A9322FAF5941DF70737CA69F152A3 ; wire I9625E96E33563830A2A0ED7263124B10 ; wire I1B43D1CE930FCA067FA31726F2C15FEE ;
wire [31:0] I697639B04C0F4B6F9764F8122329FB7C ; wire [IC6E51C590A86FEEF8592133ED3A689E7 - 1:0] I11AAD529B8C632E2B3F7E5810F154FAE ;
wire [I9A19F862D1FD27BAC93F9AC85F8F1B2B - 1:0] I6E8F4533B895189C22AD2D5F06D2C022 ; wire [IB985C42C0963EF96E8DAFEE1BF657C01
- 1:0] IB9BCD6E1EA621FDF5DD229996ADC5F8F ; wire [I8224701A907960C6458368B9E178E270 - 1:0] I6037B76B56AF44132A3D98CA48DE55B0 ;
wire [gx_ipx_data_sz - 1:0] I9A5D7FA3649743F4C12D7A2A0F5D00B9 ; wire IB72EDE3F33BC320C4BB54A891CA0124E ; wire I597BFE708F080A1AC7F68B18B2D32AEF ;
wire I452B7C3155C15AA425E22E8ACF0B4BDF ; wire IBCEC5B979CD682F2C507E946AAC6F86F ; wire I443AE8A2A80F3D4BC5B0F9739DC268B7 ;
wire IF35D2DA8FDBB83C8C227111A766BE7D7 ; wire I026F76BAC2C8DF5D427631DEA76B062F ; wire IE9523C108AFE8D1C07903BFCE449B9F8 ;
wire IFD9B46ACBF1F17D2A8C784B3B4B2901E ; wire I42C3C6068A9CD9CB33558F95CD336652 ; wire I39F7612EB75C5A11AF508BF344CD51B8 ;
wire ICF4A96ABEB44A00DC9123A0C152DC218 ; wire [IB18B8E96B09D7E54E97338C01ECBF348 - 1:0] I6C86D46877E4F106568E7404A48B3614 ;
wire [1:0] I1EBAB68345C1F3BB0BA0E7EF6A0A1648 ; wire [2:0] I25EB4135E1552B388D1686480F82F884 ; wire [gx_nr_wb_tgts
- 1: 0] IECA17FE57E485E6400F2DB42821DD251 ; wire [31:0] I02736097A9414A8EE96C59AC2C4D85D6 ; wire [3:0] IE7216A06BFCE79862D756B0F69D722FB ;
wire I109964893AEF92F63170615855D13B10 ; wire I2407989C7097E49E194FF778C1BA69FD ; wire IFDE36B1D5ECEDDC8E1D64BAC3AB778F5 ;
wire [gx_wbm_data_sz - 1:0] IF61A4C9125864F891B9412F7F8A38722 ; wire [7:0] IFDD7175F3E1142C3A73A9731A4DF519B ; wire
ICCEE7A1D3C2702A0766B02D0E4CD1F5A ; wire IF35E88F0598148E05EAD3AB0F7ED2F9E ; wire I7A68BADCCB87652618C1488B18D4A938 ;
wire [gx_wbs_data_sz - 1:0] IE5A769A04E820A9426CF9BB3B0A13E3C ; wire I5257580F4980618A2A58EA7899EEC7B5 ; wire ICBA9D9788BB5A0277607D0E038FE4333 ;
wire [gx_wbs_data_sz - 1:0] I10A77B5F026A0F0CC0D1B6C8CD9C0746 ; wire ID0B88392A9310E618D259D3AE74555DF ; wire IAB567E212EF35BD2AA033B83F2307D63 ;
wire [gx_wbs_data_sz - 1:0] IC3E05B0E9AC8F202F65F1764031827B8 ; wire I25B75CE7CA22EBCC6B686F9FD442035C ; wire IADAF74E73FA3BF461BB558E703D7C71C ;
wire [gx_wbm_data_sz - 1:0] I81A897F1890AB384489CA6655F3A90F9 ; wire I5EB48F61C7554EB021FC36EC1077B4B1 ;  assign
ox_dec_adr = I220A96CF74656D5120C8D113E4B1ED55 ; assign ox_dec_bar_hit = {I31980ABC07D19BA89784085C7754DE42 , IB55475954FE95F83F22B1C2FB76FAEC7 ,
I5078F81AE0F5DCD4CC2ABEE2CEF9C827 , IF9A16909C25386742335A246DEDE12E8 , IFFF50035216FD68A74F8164F0EE74689 , IA6774F4F4F3AF83C6A9E233DB00F89A0 };
assign ox_dec_func_hit = IE1F9397E899B4E938A0D54FC51445C13 ; assign ox_ipx_cc_npd_num = IF60FDFFF213C716383F950A9422A1758 ;
assign ox_ipx_cc_pd_num = I4FF065235743696A883B835CA5B1B85D ; assign ox_ipx_cc_processed_npd = IA4F8AA6824642C6A9DC9A7747287580D ;
assign ox_ipx_cc_processed_nph = I010A8CBEA176E0F2178CBA8B77E6FE07 ; assign ox_ipx_cc_processed_pd = I00B00319AA148C3D5F9C641ABDDBAFA3 ;
assign ox_ipx_cc_processed_ph = I92625F81A8AD6C4657526FD7E7F0D00C ; assign ox_ipx_tx_data = I9A5D7FA3649743F4C12D7A2A0F5D00B9 ;
assign ox_ipx_tx_dwen = IB72EDE3F33BC320C4BB54A891CA0124E ; assign ox_ipx_tx_end = I597BFE708F080A1AC7F68B18B2D32AEF ;
assign ox_ipx_tx_req = I452B7C3155C15AA425E22E8ACF0B4BDF ; assign ox_ipx_tx_st = IBCEC5B979CD682F2C507E946AAC6F86F ;
assign ox_wbm_adr = I6C86D46877E4F106568E7404A48B3614 ; assign ox_wbm_bte = I1EBAB68345C1F3BB0BA0E7EF6A0A1648 ;
assign ox_wbm_cti = I25EB4135E1552B388D1686480F82F884 ; assign ox_wbm_cyc = IECA17FE57E485E6400F2DB42821DD251 ;
assign ox_wbm_dat = I02736097A9414A8EE96C59AC2C4D85D6 ; assign ox_wbm_sel = IE7216A06BFCE79862D756B0F69D722FB ;
assign ox_wbm_stb = I109964893AEF92F63170615855D13B10 ; assign ox_wbm_we = I2407989C7097E49E194FF778C1BA69FD ; assign
ox_wbs_ack = IAB567E212EF35BD2AA033B83F2307D63 ; assign ox_wbs_dat = IC3E05B0E9AC8F202F65F1764031827B8 ; assign
ox_wbs_err = 1'b0; assign ox_sys_rst_n = ID872B1CCC580E5915A782E136C7A691B ; assign ox_sys_rst_func_n = ~IB1AAAED8469CADFA3AB4BF806A8466B6 ;
 assign I25B75CE7CA22EBCC6B686F9FD442035C = I09D474E43198BB26D683E473E35C90C8 & IA51154D40B341A92D3FF48956FE47EDD ;
assign IADAF74E73FA3BF461BB558E703D7C71C = IFDE36B1D5ECEDDC8E1D64BAC3AB778F5 | I1B43D1CE930FCA067FA31726F2C15FEE ;
assign I81A897F1890AB384489CA6655F3A90F9 = IF61A4C9125864F891B9412F7F8A38722 | I697639B04C0F4B6F9764F8122329FB7C ;
assign I5EB48F61C7554EB021FC36EC1077B4B1 = IB6F57A3FE1F5B6A182168AC92AC3D457 & (|IDCB78AD56EF8FEF35AAF4DED8D1F87B6 );
 IA68D2B0762B11205E05F2AB6538CBB65 #( .IB71844FFA3AB85FEF45EAB4D35395752 (IB89F6B40906A7C6F23E0C9CD1176DAD6 ), .IDB751C3DD512B8355CF27001F983880A
(gx_ipx_data_sz ), .I66C185998F46A7148163982E39BCD296 (gx_tech_lib ), .IE33DC83D2AA8913B2CB48378DAF2547A (gx_wbm_data_sz )
) IB07EBEEDDFB2F1AD47B27590E82A92BE ( .ICCFB0F435B37370076102F325BC08D20 (ix_clk_125 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(ix_rst_n ), .I93AE636CE82DE94CB11ACCF59F8C2254 (ix_ipx_dl_up ), .I2AED852F071D7FF5A04BEFAF4E7F3B0F (ix_ipx_rx_data ),
.I9B9FF20B523F68871F4D27848F9B4E44 (ix_ipx_rx_end ), .I694FF88E6CB22CE905A2A9A9E00AF7F1 (ix_ipx_rx_st ), .ID637623B1855D5BBD98CB5D56E107619
(IAF786EDCB7BC54665688D1FC2E0E922F ), .IA05976160EBA6DEFAAAA66970A81B32D (IB552918C70C5F8374FC906E0C2225F89 ), .IF249B786312150CAA567D0B3F1DC760E
(IE593D61A89622FBF1D4D61DBF77B0759 ), .I99A7C01D853D4CD1BF86EA17B055AE82 (IEB0657AD1CF8431866F1DACFA91DAE9C ), .IAB7D8322CEA20D7B2FC0EF19A061CB19
(I09D474E43198BB26D683E473E35C90C8 ), .I14B85FB28FCEF458E6F9665F2960F9A2 (IA51154D40B341A92D3FF48956FE47EDD ), .I5F4B958B42F630F4DF0F2B5578E72A4C
(I2FB68C8CAC3EE2BC47F461C034FBC722 ), .I08C693C25A115282C35BE10561F37009 (I78FE781BC8B5C49E9E0559250B6D4289 ), .ID7A2A8B1E9D92B60194D5FAFAAB15208
(IA5B0FE243F631FAA054C108CC3F72E10 ), .IFAF3E1E717F33D0636699473D114FAAC (IE228EF2D803387145092976501986E10 ), .I89CFFA73C7546481B72B0FB06D799AEE
(I6DF8AFD2D5E8EFB85D4507AC54B8E25C ), .I3E859D8CBD08E747693AC2BA98F2B947 () ); generate if (gx_wbm_data_sz == 32)
begin : IBC36250DA2BF94F52180778260423E0E I4CACC63B64035D749DE3C4BCF79F626C #( .IA0709F456132ABB4EB324E1598AAB825
(IB89F6B40906A7C6F23E0C9CD1176DAD6 ), .IFC796EA7F9507A2288E499F7B9ECC63E (I90D984439DDA58639C67AC709C0E6CC9 * I249BB13F12A1B213E14013F118AB1013 ),
.IDB9D60794264C5F8E5363941194A797B (gx_nr_wb_tgts ), .I50AC25E9687F891BB7188EED025C1323 (I37BDD1A019498B0050A3FF971DCE0165 ),
.ID7C7F9F2E39BEBEE2ACFA8040034E48D (IB18B8E96B09D7E54E97338C01ECBF348 ) ) I94FE2407114DC63C56410ECFC239E4D4 ( .ICCFB0F435B37370076102F325BC08D20
(ix_clk_125 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7 (ix_rst_n ), .I69B8FD7561F9CA8AAF4E50C5B2DCF850 (IFD9B46ACBF1F17D2A8C784B3B4B2901E ),
.IA85D446CD214F6B3CE6418205432D870 (I42C3C6068A9CD9CB33558F95CD336652 ), .IBB8FE5B389C0BD7BA64F2E05FCDC4485 (I39F7612EB75C5A11AF508BF344CD51B8 ),
.I45A8F29589769D54C9D702481065CB45 (ICF4A96ABEB44A00DC9123A0C152DC218 ), .IFF5E23C5A17BB678C108274E28C56424 (I395C5996AD91572D0F6652373B6018E7 ),
.IDE425A12275C43D9056DCF647A2D8258 (I5B507E107F91FDBF0B2EEF7DD9AE40C5 ), .I65B14714ECFCC218D3A788DF7696216B (IBAE868C7DE15BF2F751B0177B798BDCD ),
.IA1F0CBEC8E9EAD83D0098DD96A1EFC32 (3'b000), .IFC18758E8987A9913FD94A5DFEE774E2 (1'b0), .IF5E7E4E58741BF3FE58442AB377ED57F
(IC0197882115D001485B37646159E234E ), .IF5B4924BEAEA6935367AC2739021882F (1'b0), .I7985A5A43CBBBC8E0D3FCFEE38DDF221
(1'b0), .I7E600D684E83043922C1FE27CC6213E4 (ix_dec_wb_cyc ), .I93AE636CE82DE94CB11ACCF59F8C2254 (ix_ipx_dl_up ),
.I9119CE851F731CBC5834D0370CCA6908 (I1BAAE01807D45E9F21D2ACB2BCB4F621 ), .I9F3623AEB414A15CECD2A8FD8791C79D (I2FB68C8CAC3EE2BC47F461C034FBC722 ),
.I36824F33FF142FDE2AFE9BC4759DB690 (I78FE781BC8B5C49E9E0559250B6D4289 ), .I5E84ED10AD623502BC750C5E797D1428 (IA5B0FE243F631FAA054C108CC3F72E10 ),
.IA886199C0F7609B072DAE171DFC98CD8 (IE228EF2D803387145092976501986E10 ), .IA067043029572C8598E352E0A66EA337 (I6DF8AFD2D5E8EFB85D4507AC54B8E25C ),
.ICB518A59CAE27DDB6398AB22F5D74259 (I11AAD529B8C632E2B3F7E5810F154FAE ), .I9F4F7E2C4A4A8FB2780021EDF6E4ADEF (I443AE8A2A80F3D4BC5B0F9739DC268B7 ),
.I07B0EBE8FBC21BDBE894D73C90EDC5AB (IADAF74E73FA3BF461BB558E703D7C71C ), .I44B3CB0FFE4214C92C98CD6ECFC52D5A (|IECA17FE57E485E6400F2DB42821DD251 ),
.I3D6C771D05CA1A769E61302C086494B8 (I81A897F1890AB384489CA6655F3A90F9 ), .IC2E260CA356C994048CCB108C7E359D1 (IF60FDFFF213C716383F950A9422A1758 ),
.IE707B5D4A74BA1BD745B52E0C07932C0 (I4FF065235743696A883B835CA5B1B85D ), .I6E70C748D9C56227AB1182F36658AE5C (IA4F8AA6824642C6A9DC9A7747287580D ),
.I59B23598E8ADE1982F184EF67BEB0979 (I010A8CBEA176E0F2178CBA8B77E6FE07 ), .I33E409903692F5ECA2EC3553F9D1659E (I00B00319AA148C3D5F9C641ABDDBAFA3 ),
.I437E57D42FB91B674CCBCC915BF9D653 (I92625F81A8AD6C4657526FD7E7F0D00C ), .I55AFDDE17B53D7F65849D39B02B07417 (),
.I65FE2DB4E1CB5A488A45D60041AB5F64 (), .I0C796C206FE7060B578156D0110461EB (I220A96CF74656D5120C8D113E4B1ED55 ),
.IFC86A6522A8CA080A0DB7F384D9CE6FA ( ), .I484F77D7967D25736EB27A0ED76CCB5F (IBE8D7D536CBDF087E7E00B93DA215E3D ),
.I7E0431D7F1A92C0ED1F030F36BF809B7 ( ), .I3E6965EC606FD6C2871F2C0993204C57 (I4DC446D96F0774A667A70D52D9392874 ),
.IFF25B820DFD457D71B32B130ABE5DA3F (I3FF9BAFBF91288E78D7EA6DD95DB3A40 ), .I20FA57C9A87CB2AA26088D9FA1743F70 ( ),
.I51C881E8B9B36D7A724BC7B8EC533957 ( ), .ID3E7F4B58943229FEE6313A36B3F8693 (IE67E5659AC07E2D371890CDACFA6ED42 ),
.I1FDEC1735547330C00A0B8DFE1FB10C3 (I18137FEBF7FA4CE04FDE793386121F57 ), .IBD6A65D48B4A68CA0D2A82F79053757B (I0B37325C0AB5EEA3148286371EB202D1 ),
.I15EC78E3DE1101BFF2B227962683E113 (IAF786EDCB7BC54665688D1FC2E0E922F ), .I7C4DADE2C05F6DCECCAF7AD6F7BF2FF8 (I6609F40DB9BF2AAD262974646AD5EBE5 ),
.IEEFA85D6664F09687B5CA591C701DC34 (IAE96F702FDFFAF4D7DD2303A7E5CAA82 ), .ID4A284C76C6EABEEBA8E0AE18003FBAC (I314F20E260B367A911975FFD9E094426 ),
.I6010C20131B976554A498745FEEEB580 (I4A399AD6EACAD372F1F0ED553AF29E10 ), .I46E8CA15DC1E8B3B2200999A53029704 (IE81C89DB2F6C737F2D82BE35AFC7DDA2 ),
.IEC45B60C7D1A49FFA84D3F5D121A2579 (IC13572948B0A4216A965E35100DE669F ), .I9AF46E2AA924FA7E0F5D7290324BABF9 (I599F86FA1B9AEED5B32EE8B27DFFFACE ),
.I59D9A9A677978229C1F87AA1A3A0C304 (I291FF0AF6B998FB4D8BD958CFDA1CF8C ), .I9301CE4E9B877D08EDBD1584D6BE017A ( ),
.I51698892CBD372EE66AF3EA4D0ECE23F ( ), .I1347408C9E757F34EA4D78F53447BD9B ( ), .I2BE88607F3C31B47400F3A35E08B7EAD
(IDCB78AD56EF8FEF35AAF4DED8D1F87B6 ), .I7D901091F9E0741061C75B54467D48A0 (IEC017B3AB9F16AE871D5253A5257D941 ), .I40EF39BB4F4F4A031C8FD1026EF53063
(I87343FD56CEFDCB10F9A272CF1F0CA8E ), .I42427E866FF31BC28E35C71EC172E26B (IB8F3718FAD7719FD71FDE3B0DE8D7445 ), .I7AEBDB3D2CD4891A528BA81F5F54B20D
(IB6F57A3FE1F5B6A182168AC92AC3D457 ), .ID16819FEAA95700005E383E7DA0C8E13 (I7681E0E609A03559F13166ACF7852905 ), .IE0337CA803FBA20F38A0CD2A900C6534
(I507A0A1A3C69E79845F5C15AFFAF6595 ), .I592A6A3BA99B09C24695C7A609F9053F (IDB0B420EA96A60B402FECD3AE3620DCC ), .I368749E68EAF9F462385FAD36180A9FE
(I678B3227DE7FFEFE726CE68123B91F8D ) ); end endgenerate generate if (gx_wbm_data_sz == 64) begin : I6A9FBF362205F11DF0825B6130C9BDE7
I1F8444FEC9FE4C651C698EE6099B529D #( .IB71844FFA3AB85FEF45EAB4D35395752 (IB89F6B40906A7C6F23E0C9CD1176DAD6 ), .IDB9D60794264C5F8E5363941194A797B
(gx_nr_wb_tgts ), .ID7C7F9F2E39BEBEE2ACFA8040034E48D (IB18B8E96B09D7E54E97338C01ECBF348 ) ) I94FE2407114DC63C56410ECFC239E4D4
( .ICCFB0F435B37370076102F325BC08D20 (ix_clk_125 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7 (ix_rst_n ), .I69B8FD7561F9CA8AAF4E50C5B2DCF850
(IFD9B46ACBF1F17D2A8C784B3B4B2901E ), .IA85D446CD214F6B3CE6418205432D870 (I42C3C6068A9CD9CB33558F95CD336652 ), .IBB8FE5B389C0BD7BA64F2E05FCDC4485
(I39F7612EB75C5A11AF508BF344CD51B8 ), .I45A8F29589769D54C9D702481065CB45 (ICF4A96ABEB44A00DC9123A0C152DC218 ), .IFF5E23C5A17BB678C108274E28C56424
(I395C5996AD91572D0F6652373B6018E7 ), .IDE425A12275C43D9056DCF647A2D8258 (I5B507E107F91FDBF0B2EEF7DD9AE40C5 ), .I65B14714ECFCC218D3A788DF7696216B
(IBAE868C7DE15BF2F751B0177B798BDCD ), .IA1F0CBEC8E9EAD83D0098DD96A1EFC32 (3'b000), .IFC18758E8987A9913FD94A5DFEE774E2
(1'b0), .IF5E7E4E58741BF3FE58442AB377ED57F (IC0197882115D001485B37646159E234E ), .IF5B4924BEAEA6935367AC2739021882F
(1'b0), .I7985A5A43CBBBC8E0D3FCFEE38DDF221 (1'b0), .I7E600D684E83043922C1FE27CC6213E4 (ix_dec_wb_cyc ), .I93AE636CE82DE94CB11ACCF59F8C2254
(ix_ipx_dl_up ), .I9119CE851F731CBC5834D0370CCA6908 (I1BAAE01807D45E9F21D2ACB2BCB4F621 ), .I9F3623AEB414A15CECD2A8FD8791C79D
(I2FB68C8CAC3EE2BC47F461C034FBC722 ), .I36824F33FF142FDE2AFE9BC4759DB690 (I78FE781BC8B5C49E9E0559250B6D4289 ), .I5E84ED10AD623502BC750C5E797D1428
(IA5B0FE243F631FAA054C108CC3F72E10 ), .IA886199C0F7609B072DAE171DFC98CD8 (IE228EF2D803387145092976501986E10 ), .IA067043029572C8598E352E0A66EA337
(I6DF8AFD2D5E8EFB85D4507AC54B8E25C ), .ICB518A59CAE27DDB6398AB22F5D74259 (I11AAD529B8C632E2B3F7E5810F154FAE ), .I9F4F7E2C4A4A8FB2780021EDF6E4ADEF
(I443AE8A2A80F3D4BC5B0F9739DC268B7 ), .I07B0EBE8FBC21BDBE894D73C90EDC5AB (IADAF74E73FA3BF461BB558E703D7C71C ), .I44B3CB0FFE4214C92C98CD6ECFC52D5A
(|IECA17FE57E485E6400F2DB42821DD251 ), .I3D6C771D05CA1A769E61302C086494B8 (I81A897F1890AB384489CA6655F3A90F9 ),
.IC2E260CA356C994048CCB108C7E359D1 (IF60FDFFF213C716383F950A9422A1758 ), .IE707B5D4A74BA1BD745B52E0C07932C0 (I4FF065235743696A883B835CA5B1B85D ),
.I6E70C748D9C56227AB1182F36658AE5C (IA4F8AA6824642C6A9DC9A7747287580D ), .I59B23598E8ADE1982F184EF67BEB0979 (I010A8CBEA176E0F2178CBA8B77E6FE07 ),
.I33E409903692F5ECA2EC3553F9D1659E (I00B00319AA148C3D5F9C641ABDDBAFA3 ), .I437E57D42FB91B674CCBCC915BF9D653 (I92625F81A8AD6C4657526FD7E7F0D00C ),
.I55AFDDE17B53D7F65849D39B02B07417 (), .I65FE2DB4E1CB5A488A45D60041AB5F64 (), .I0C796C206FE7060B578156D0110461EB
(I220A96CF74656D5120C8D113E4B1ED55 ), .IFC86A6522A8CA080A0DB7F384D9CE6FA ( ), .I484F77D7967D25736EB27A0ED76CCB5F
(IBE8D7D536CBDF087E7E00B93DA215E3D ), .I7E0431D7F1A92C0ED1F030F36BF809B7 ( ), .I3E6965EC606FD6C2871F2C0993204C57
(I4DC446D96F0774A667A70D52D9392874 ), .IFF25B820DFD457D71B32B130ABE5DA3F (I3FF9BAFBF91288E78D7EA6DD95DB3A40 ), .I20FA57C9A87CB2AA26088D9FA1743F70
( ), .I51C881E8B9B36D7A724BC7B8EC533957 ( ), .ID3E7F4B58943229FEE6313A36B3F8693 (IE67E5659AC07E2D371890CDACFA6ED42 ),
.I1FDEC1735547330C00A0B8DFE1FB10C3 (I18137FEBF7FA4CE04FDE793386121F57 ), .IBD6A65D48B4A68CA0D2A82F79053757B (I0B37325C0AB5EEA3148286371EB202D1 ),
.I15EC78E3DE1101BFF2B227962683E113 (IAF786EDCB7BC54665688D1FC2E0E922F ), .I7C4DADE2C05F6DCECCAF7AD6F7BF2FF8 (I6609F40DB9BF2AAD262974646AD5EBE5 ),
.IEEFA85D6664F09687B5CA591C701DC34 (IAE96F702FDFFAF4D7DD2303A7E5CAA82 ), .ID4A284C76C6EABEEBA8E0AE18003FBAC (I314F20E260B367A911975FFD9E094426 ),
.I6010C20131B976554A498745FEEEB580 (I4A399AD6EACAD372F1F0ED553AF29E10 ), .I46E8CA15DC1E8B3B2200999A53029704 (IE81C89DB2F6C737F2D82BE35AFC7DDA2 ),
.IEC45B60C7D1A49FFA84D3F5D121A2579 (IC13572948B0A4216A965E35100DE669F ), .I9AF46E2AA924FA7E0F5D7290324BABF9 (I599F86FA1B9AEED5B32EE8B27DFFFACE ),
.I59D9A9A677978229C1F87AA1A3A0C304 (I291FF0AF6B998FB4D8BD958CFDA1CF8C ), .I9301CE4E9B877D08EDBD1584D6BE017A ( ),
.I51698892CBD372EE66AF3EA4D0ECE23F ( ), .I1347408C9E757F34EA4D78F53447BD9B ( ), .I2BE88607F3C31B47400F3A35E08B7EAD
(IDCB78AD56EF8FEF35AAF4DED8D1F87B6 ), .I7D901091F9E0741061C75B54467D48A0 (IEC017B3AB9F16AE871D5253A5257D941 ), .I40EF39BB4F4F4A031C8FD1026EF53063
(I87343FD56CEFDCB10F9A272CF1F0CA8E ), .I42427E866FF31BC28E35C71EC172E26B (IB8F3718FAD7719FD71FDE3B0DE8D7445 ), .I7AEBDB3D2CD4891A528BA81F5F54B20D
(IB6F57A3FE1F5B6A182168AC92AC3D457 ), .ID16819FEAA95700005E383E7DA0C8E13 (I7681E0E609A03559F13166ACF7852905 ), .IE0337CA803FBA20F38A0CD2A900C6534
(I507A0A1A3C69E79845F5C15AFFAF6595 ), .I592A6A3BA99B09C24695C7A609F9053F (IDB0B420EA96A60B402FECD3AE3620DCC ), .I368749E68EAF9F462385FAD36180A9FE
(I678B3227DE7FFEFE726CE68123B91F8D ) ); end endgenerate IAC6C4C771C836211892F0FD3F47BC076 #( .I857673E5DE2CF777499EE369473CBCCC
(gx_cs_f0_bar0_size ), .IA874AED52F9C16F13B580898DA0E85AC (gx_cs_f0_bar0_is_64_bit ), .I45E74A319CD545DA84EE876844F12DF8
(gx_cs_f0_bar0_is_io_space ), .I212658651766EFCF73257AF1E3121AF8 (gx_cs_f0_bar0_is_prefetchable ), .I2610FF174BEEE098C8D9C9374191F122
(gx_cs_f0_bar1_size ), .IA8729443C3DAFAFDD37A6BED4B24F26C (gx_cs_f0_bar1_is_io_space ), .I08EC85B0527EBF111FDA96E4BD71B6BF
(gx_cs_f0_bar1_is_prefetchable ), .I6C75B7796A1597A63620710B69C04958 (gx_cs_f0_bar2_size ), .I86AD8EB6B8FA8A1AA6EA64DE4357E4EA
(gx_cs_f0_bar2_is_64_bit ), .I5C0FF6EA47D5544D48B9200C35F2015D (gx_cs_f0_bar2_is_io_space ), .IED6EFA8FE915B71B8E198535343CFBFB
(gx_cs_f0_bar2_is_prefetchable ), .I98F26EACDFB5625667BCAFBDB2867748 (gx_cs_f0_bar3_size ), .I3CAEAE4A6B7BA30F88F0945373893582
(gx_cs_f0_bar3_is_io_space ), .ICC1064DA289312A92936196EA26F0023 (gx_cs_f0_bar3_is_prefetchable ), .I78F9B7090517BBEEBC1543199FBA4D34
(gx_cs_f0_bar4_size ), .I731C578B2B8A6173399D3CABA7E98889 (gx_cs_f0_bar4_is_64_bit ), .IE18DEDE16538C154B2EFCB2652C25FD5
(gx_cs_f0_bar4_is_io_space ), .IB6EB169241E23C32C11DDDC27322BCE6 (gx_cs_f0_bar4_is_prefetchable ), .I83476C8D11033DBF952882C55FC0E55B
(gx_cs_f0_bar5_size ), .I156838D82D20DC7C269685B24CB4A8B0 (gx_cs_f0_bar5_is_io_space ), .I86134D1B828E3E59B9C4B66EC0920D98
(gx_cs_f0_bar5_is_prefetchable ), .IC2EB58967FBD1CD5C54491738F4BAD86 (gx_cs_f0_class_code ), .IBBBF11BAEEC8458B08DFB6E2D9D1C850
(gx_cs_f0_device_id ), .IA54DA90446D375855AF33292D2570A3C (gx_cs_f0_int_count ), .IAD54DD4DF3ABBB4563A2B75498325CD7
(gx_cs_f0_int_pin ), .I02756A8C58D5B37B7049B7F6FA2073B7 (gx_cs_f0_revision_id ), .I1066D287D755AADD24EE379E400F8DA8
(gx_cs_f0_subsystem_id ), .IE8C1215A45516D3178A8A93152E05EE2 (gx_cs_f1_bar0_size ), .I6A67F4FE467D33BBE90E5158D72171A4
(gx_cs_f1_bar0_is_64_bit ), .I8F998DCDBE9627EA583F7BB408EC780D (gx_cs_f1_bar0_is_io_space ), .I8695C513BA5D9DA307CC481D6AFFB133
(gx_cs_f1_bar0_is_prefetchable ), .IEE21CD471C5E4E6CE83A164513BC7722 (gx_cs_f1_bar1_size ), .I56DA37D670BDECB81356B81560DC8649
(gx_cs_f1_bar1_is_io_space ), .IB36C0E6BB9CF8D4E4A2F31086369A6EC (gx_cs_f1_bar1_is_prefetchable ), .I6C4BB963A9FEECAA07E250007DE29E69
(gx_cs_f1_bar2_size ), .I7725F462040C54BFDFC296100F95D5D0 (gx_cs_f1_bar2_is_64_bit ), .IC022347DC0BBA44450EA061654CE4130
(gx_cs_f1_bar2_is_io_space ), .I8DFF460C39C720D8E01DF9AD54E62457 (gx_cs_f1_bar2_is_prefetchable ), .I128970AF889EC52F4195C246A49524BA
(gx_cs_f1_bar3_size ), .I61E4D6D4FFCCB1C283902514C76CD3AA (gx_cs_f1_bar3_is_io_space ), .ID0832173F4D69F0B96DB00FA9805F75F
(gx_cs_f1_bar3_is_prefetchable ), .I171E938E7CDE23987F02EB923184A5C3 (gx_cs_f1_bar4_size ), .I5A509B803B47567D6FA4F4CB4C6AA95D
(gx_cs_f1_bar4_is_64_bit ), .I2C1FDD71B618A0C398964466A5958BF0 (gx_cs_f1_bar4_is_io_space ), .ICE7C691E1DC04B92371B76DCE234C732
(gx_cs_f1_bar4_is_prefetchable ), .IA9D9F2D7EEC92A228D6CC71EE9A86E0E (gx_cs_f1_bar5_size ), .I7356A0718B40AEF099CE99273A8CBC19
(gx_cs_f1_bar5_is_io_space ), .I4521B8E3C71C6E5D7639756B81D56C58 (gx_cs_f1_bar5_is_prefetchable ), .IB52E64F4A5E8239ED2BF949AC0702ACE
(gx_cs_f1_class_code ), .IA5A53C930B674A8F9761966972CFB6F6 (gx_cs_f1_device_id ), .I97F18A3381F2546EB21E07DF7628912F
(gx_cs_f1_int_count ), .I2FCDB5B825200EDE4D7757A0621663E0 (gx_cs_f1_int_pin ), .IE50492CEE03959C13AD5E521CC7F2FEF
(gx_cs_f1_present ), .IC745524098FFC5FBA778DA59D2444D9B (gx_cs_f1_revision_id ), .I7507C2B666C444A66EDA2CFDB6DCEEB9
(gx_cs_f1_subsystem_id ), .I1A39FC80F18CFB225DD25F1158A43FEB (gx_cs_f2_bar0_size ), .IFA1CC1A50C8D64B9481E806D15AF3CA5
(gx_cs_f2_bar0_is_64_bit ), .IF089B8BB6C2663DE1CA53AB4AB67231B (gx_cs_f2_bar0_is_io_space ), .I348F387B0CC3540AF0215535F676D5A2
(gx_cs_f2_bar0_is_prefetchable ), .I3AB6DCBD252A38D5954C33DB9CFA020B (gx_cs_f2_bar1_size ), .IFE55C92252D5A4FCF3878CC98FCAD612
(gx_cs_f2_bar1_is_io_space ), .IC2181A40E4750EEA118AA81ABB4E415B (gx_cs_f2_bar1_is_prefetchable ), .I813CE6D8049DC9123C58691D1DA81B59
(gx_cs_f2_bar2_size ), .I50243AFBCB64F92A3F6EEC157034F4FC (gx_cs_f2_bar2_is_64_bit ), .I38E6C6DF2535A2049746702855108B5A
(gx_cs_f2_bar2_is_io_space ), .I0FFEAFBF23F15260885D040F12B66960 (gx_cs_f2_bar2_is_prefetchable ), .I31E80F0EE05B52A92941F617BDCEF890
(gx_cs_f2_bar3_size ), .I509611AF740C942BA82FB9ECE7BA4E67 (gx_cs_f2_bar3_is_io_space ), .I586C95E6CCC79680B179527AE8977C4E
(gx_cs_f2_bar3_is_prefetchable ), .I39D41D0CFF63339D485BDBCDBC3A8729 (gx_cs_f2_bar4_size ), .IF833CBC3D7A215E6C5635F3F07A09365
(gx_cs_f2_bar4_is_64_bit ), .IE106099B16008BAE163236DC5CF4EAFE (gx_cs_f2_bar4_is_io_space ), .IC4C3CD51A29DC2F222334D23407BB4E7
(gx_cs_f2_bar4_is_prefetchable ), .I7C988FF99F8B28AB1CE2299774306236 (gx_cs_f2_bar5_size ), .I4FF1FE282379DCB83A2AF4F7A12AF6CA
(gx_cs_f2_bar5_is_io_space ), .IB5B3486ECA0F911FF5D92A37ECF53B4A (gx_cs_f2_bar5_is_prefetchable ), .I0B5E80731173820DE30A1D6C548B918B
(gx_cs_f2_class_code ), .I8A848F283F0A33BC04B5173E5E3FE015 (gx_cs_f2_device_id ), .I0069A39965C0330678D64B612F60F78D
(gx_cs_f2_int_count ), .I30A298A8327798F01C20DDAD6A556FB3 (gx_cs_f2_int_pin ), .I0B3C14F69FAC563649E26679A3D8B1CD
(gx_cs_f2_present ), .I4EB1044CFC38A54424DBAA59B9641ED6 (gx_cs_f2_revision_id ), .IC920957C9C4BA12361B2EB75CD52EA74
(gx_cs_f2_subsystem_id ), .IB231E22D146559D11318B25AE0BA8C7A (gx_cs_f3_bar0_size ), .I7377F8B5325C7EE7D12D8B4B6A18183F
(gx_cs_f3_bar0_is_64_bit ), .I17C1305CE886D24D942A2A62C4DB3617 (gx_cs_f3_bar0_is_io_space ), .ID926607BDA4008824BC8A9A1B67C04B7
(gx_cs_f3_bar0_is_prefetchable ), .IE4511A2FC6AD3FBAEAADD1EF75F0B773 (gx_cs_f3_bar1_size ), .I0B29563399BE9E04B2FE3DE714C7DCE6
(gx_cs_f3_bar1_is_io_space ), .I698853A251199BE8A5753717E876DA52 (gx_cs_f3_bar1_is_prefetchable ), .IA3BC4D015F529FD7E88E1370A882D0DF
(gx_cs_f3_bar2_size ), .I3463AC2A02018CF2288043A9C3E47A4F (gx_cs_f3_bar2_is_64_bit ), .IFDC235A84B81F7EB6EA5B1ED1F71197F
(gx_cs_f3_bar2_is_io_space ), .IF0C0D849F42A4C05A7BF373811D5F5F5 (gx_cs_f3_bar2_is_prefetchable ), .I59B19D300B55C10DB1B10364E9E59201
(gx_cs_f3_bar3_size ), .IB1CD9FD007D322042A1087AC76B782B4 (gx_cs_f3_bar3_is_io_space ), .I6A959CC2CFE148A0D8579A1CEE0C6699
(gx_cs_f3_bar3_is_prefetchable ), .I1953E43D30396B1EDBD48DAD13C6A240 (gx_cs_f3_bar4_size ), .IC02B62ACA36F1FEBB031FE435BA48A9A
(gx_cs_f3_bar4_is_64_bit ), .IAE6C36DBDB6FF8E962D96D8F1FB95CC1 (gx_cs_f3_bar4_is_io_space ), .I82E91D4ACF151209B3234E6F867049F1
(gx_cs_f3_bar4_is_prefetchable ), .I9806BFEA675277E4572CB4FD0C9C0D8C (gx_cs_f3_bar5_size ), .I802B81175874E1E34C3E4EE6C7F0B969
(gx_cs_f3_bar5_is_io_space ), .I00773A8B25BA28541FF04BC530185E7F (gx_cs_f3_bar5_is_prefetchable ), .IB2267C4E34709B9CE9D697340B9DA12F
(gx_cs_f3_class_code ), .I37AC0331E13434E399C90A5408FB09E2 (gx_cs_f3_device_id ), .IC69BEB80DB094A65F3DFB0265F8616DE
(gx_cs_f3_int_count ), .I6C4A37BD8E4A0A1D9639A3FA64D5F8C3 (gx_cs_f3_int_pin ), .IFA272F301A5935EE15CB134524665363
(gx_cs_f3_present ), .ID969B30E2BD8213873A2D19FFDEF204A (gx_cs_f3_revision_id ), .IC3F1AF003F5E2257563771F88647B5FF
(gx_cs_f3_subsystem_id ), .I21752C34E9BF9458DB0D20BA11A8898B (gx_cs_f4_bar0_size ), .IBFD9199C154D56895B673A496CF82DA3
(gx_cs_f4_bar0_is_64_bit ), .I900E9757930519C7865CA2247E6CC23A (gx_cs_f4_bar0_is_io_space ), .IFA7D0D435AE6BBF59445626F82B8B26E
(gx_cs_f4_bar0_is_prefetchable ), .IA794CD2FEB24AB956EC1914852D2E7D5 (gx_cs_f4_bar1_size ), .IAED1399D2D60713A0101069DD427D0A0
(gx_cs_f4_bar1_is_io_space ), .I72E6ED810779933C7E2125FC345DEC0B (gx_cs_f4_bar1_is_prefetchable ), .I3C7842C10567F9851F14519598E7EE93
(gx_cs_f4_bar2_size ), .I1DE5880AD46DABF7282A3FF245F71602 (gx_cs_f4_bar2_is_64_bit ), .I7747208BC7A624CD71D5BB421E9EE4A4
(gx_cs_f4_bar2_is_io_space ), .I4103D81EBFB4946FA8F9593A8B7DE5C8 (gx_cs_f4_bar2_is_prefetchable ), .I858B464778E6994385995C3205FB37B0
(gx_cs_f4_bar3_size ), .I785E686713BEF380843045D4DB00E51C (gx_cs_f4_bar3_is_io_space ), .IABD30C53E56587015015FE5F556929D7
(gx_cs_f4_bar3_is_prefetchable ), .IABB4198D13BE4058E856EBC11D8D6565 (gx_cs_f4_bar4_size ), .I0405497FA63FB5AA449F0C813D8E8F89
(gx_cs_f4_bar4_is_64_bit ), .I6F86DD61D81AE7AE015C945BA5CF8828 (gx_cs_f4_bar4_is_io_space ), .I69C4352219E15BD98C0B6A7428BAB037
(gx_cs_f4_bar4_is_prefetchable ), .I68ED8551754B5BAA65EB2F191A697C4B (gx_cs_f4_bar5_size ), .ICE0C22941CF3ECFDB4B47576E4E4A06E
(gx_cs_f4_bar5_is_io_space ), .I262F500CDAF1182E64A895FA5F58D006 (gx_cs_f4_bar5_is_prefetchable ), .ID88F3DF54AD4CA3D33C94EC1E1B5BB01
(gx_cs_f4_class_code ), .I8F019158F18BA70FE5953E859D4BA891 (gx_cs_f4_device_id ), .I4046611EA3EEF60ACE26738C818FDBA2
(gx_cs_f4_int_count ), .I78E815C8C6F11755E08393F339C5E874 (gx_cs_f4_int_pin ), .IE690B7723F136DA02896C0728DDADB49
(gx_cs_f4_present ), .IC377F0EF36016932385B3B0988B91B0F (gx_cs_f4_revision_id ), .IBDEA2513680CC11B2E5E42FB17332F70
(gx_cs_f4_subsystem_id ), .IDC77C35F0E8480627E0F64F68D8A39ED (gx_cs_f5_bar0_size ), .I110F59F054A1064BFB27909E2370F028
(gx_cs_f5_bar0_is_64_bit ), .IED76B05540143124D123636B36A006DA (gx_cs_f5_bar0_is_io_space ), .I96B06C30CEFF410BD39B69C003D2AC2B
(gx_cs_f5_bar0_is_prefetchable ), .I2050954950618B2F390C43E2A3A4A814 (gx_cs_f5_bar1_size ), .I3F39386711BA6D94D8C7A1C5710875D6
(gx_cs_f5_bar1_is_io_space ), .I3011FF9154FC5D6F394688805C3D9B33 (gx_cs_f5_bar1_is_prefetchable ), .I08E7BC06415AD0F55BE9EFFEB79B0315
(gx_cs_f5_bar2_size ), .IB069DEA93E56D26CAB0E5B9C9E284CDE (gx_cs_f5_bar2_is_64_bit ), .I5F80A9459505144CBBE328F0713782CC
(gx_cs_f5_bar2_is_io_space ), .IC88E0007329C31C00B55FD745AAD6590 (gx_cs_f5_bar2_is_prefetchable ), .I102247373FC0AC7EA52B3EFB2A5CC280
(gx_cs_f5_bar3_size ), .I750129419895285C7D4ABEB3C2FEEE71 (gx_cs_f5_bar3_is_io_space ), .I2CFDEF4EE4DDBFD88BE646118F3E6FE2
(gx_cs_f5_bar3_is_prefetchable ), .ID42754EA33A6C985294D5AD602396DA3 (gx_cs_f5_bar4_size ), .I6FBC4AA1ED36E030778F1A24E9C9B2E4
(gx_cs_f5_bar4_is_64_bit ), .I15A258E402E001F63FAB5BE8DF569399 (gx_cs_f5_bar4_is_io_space ), .IA2FE22B25B2F0C96B10399B2FB4B7C81
(gx_cs_f5_bar4_is_prefetchable ), .I36E46FAD7B2BA4DF9270A70F4921CC43 (gx_cs_f5_bar5_size ), .I0500A389ECC6C6D86EA16632126031AD
(gx_cs_f5_bar5_is_io_space ), .IFF2CDD869828E984763A775FF1821810 (gx_cs_f5_bar5_is_prefetchable ), .I4A7FAB30233B5A9954B6B6AD08DCADAA
(gx_cs_f5_class_code ), .IC7B583F6D8F8A6C3C62D45FA87D50A19 (gx_cs_f5_device_id ), .IAE03DAE231BA40E8DD1C02D38068EF8A
(gx_cs_f5_int_count ), .IB842E33563B3EE1795267FE015C7B1A0 (gx_cs_f5_int_pin ), .I55BE27080C370AF723A4FE096014E875
(gx_cs_f5_present ), .I229F764F8E53B82969E0B6B9234098CF (gx_cs_f5_revision_id ), .IA9807BAB69B1AFAF9739BF86D99A92C3
(gx_cs_f5_subsystem_id ), .IF02D8DF664D45B9699745A4C477F4220 (gx_cs_f6_bar0_size ), .I553DE26948BD8999C232161660D3E8AF
(gx_cs_f6_bar0_is_64_bit ), .IB99020DD53AEEF55E5DA5BF15890E9A5 (gx_cs_f6_bar0_is_io_space ), .I0108C021E74AB8DE1357A170111B08CF
(gx_cs_f6_bar0_is_prefetchable ), .IDED06CF1ED1692C601F91B904599696F (gx_cs_f6_bar1_size ), .I7926E122D54A321BCD3309E19D9A0183
(gx_cs_f6_bar1_is_io_space ), .I48C74401BD4D3F04619117E263213AFA (gx_cs_f6_bar1_is_prefetchable ), .I40F4EF6A18605258D6F6893B593AA318
(gx_cs_f6_bar2_size ), .IAB56F2CB5ED41158B5A0ABE2FD915084 (gx_cs_f6_bar2_is_64_bit ), .I11F59D9A3377C9C28FB84219B4A4E4DC
(gx_cs_f6_bar2_is_io_space ), .I3BE4D977225B6255BC284FA193DD9241 (gx_cs_f6_bar2_is_prefetchable ), .I6A49481E89496C888774F840785C0BA4
(gx_cs_f6_bar3_size ), .IE19B87A06C26E07981B4C116F5E878F7 (gx_cs_f6_bar3_is_io_space ), .IF587F6E4A635FC1DA01C698D24B80510
(gx_cs_f6_bar3_is_prefetchable ), .IBF68DF087726DF134221B625725579B8 (gx_cs_f6_bar4_size ), .I9F10A6A60E1AEDF0BC22B2ED2686E4C2
(gx_cs_f6_bar4_is_64_bit ), .I10394C1F82392903C22C104CEC600C4E (gx_cs_f6_bar4_is_io_space ), .IE4A74A61CDC56044C199B3C3D606B08E
(gx_cs_f6_bar4_is_prefetchable ), .ICE73FC6522779AED50B02BB41E81D717 (gx_cs_f6_bar5_size ), .I25D595F391F999FD69AB7E7B5B1FA99C
(gx_cs_f6_bar5_is_io_space ), .IAE37CBAA4815C82EA96E8FA0802F7443 (gx_cs_f6_bar5_is_prefetchable ), .I50BD52F5094656ECEC3714E0BAE6B0DA
(gx_cs_f6_class_code ), .IC781EE34DC62D08174F1793A9E3131B5 (gx_cs_f6_device_id ), .I7568F6D9A53738CCE095CE231BAB3F85
(gx_cs_f6_int_count ), .ID23C9147B8CA6684051791F38B473984 (gx_cs_f6_int_pin ), .IB2560D175E4507798B84D6E659FD6373
(gx_cs_f6_present ), .ID873CC05798FE57AF43DD3C4E138769B (gx_cs_f6_revision_id ), .I70E83CF258ED794C3E9EDE1260BF5578
(gx_cs_f6_subsystem_id ), .IFB72ECF29D30B02049C030502F330CE7 (gx_cs_f7_bar0_size ), .I7E6B00724A48BA5DD1C5E397542EDDC2
(gx_cs_f7_bar0_is_64_bit ), .I5C146FC803FDD1163A6BAEA53E6C5468 (gx_cs_f7_bar0_is_io_space ), .IE3404D24C7B1FA263F2EACB5CC85BFF6
(gx_cs_f7_bar0_is_prefetchable ), .IB23260A86DA99A28163B5E233CA42605 (gx_cs_f7_bar1_size ), .IEF68A43ED89112E53191106DBA0EF113
(gx_cs_f7_bar1_is_io_space ), .I95CE19A3BB94C8A24A8E3F3482EF6425 (gx_cs_f7_bar1_is_prefetchable ), .I7A84A5F1499409083F731D2A584D2D42
(gx_cs_f7_bar2_size ), .I76069160333C4C8E92944FC3A3827ED6 (gx_cs_f7_bar2_is_64_bit ), .I8EF5BB87B22B910665D13A80C6724D14
(gx_cs_f7_bar2_is_io_space ), .IFA5339CE0FEDFF3B45CF3C0167564EA1 (gx_cs_f7_bar2_is_prefetchable ), .ID3A400426A266A6F4E75F7686B9028CD
(gx_cs_f7_bar3_size ), .I071A2CF414FF8A814D779E1F54247BF1 (gx_cs_f7_bar3_is_io_space ), .I3F7B58F167F56FB985F8908CA1B7E3AE
(gx_cs_f7_bar3_is_prefetchable ), .I62A26688D23065F69E9B9D6339AA01A5 (gx_cs_f7_bar4_size ), .IE4774E19FB83A84DBF540368C45EA3A3
(gx_cs_f7_bar4_is_64_bit ), .I5ACFA0E62CCC520EE4DA1BA399F1B7E6 (gx_cs_f7_bar4_is_io_space ), .IF1CB2B99D8669C68B68BC468C83323DF
(gx_cs_f7_bar4_is_prefetchable ), .I245B45EC852C565EDD1AAC06E80DABD2 (gx_cs_f7_bar5_size ), .I59DF7AA363A19A361E3A844AD6039C40
(gx_cs_f7_bar5_is_io_space ), .IAF2433492FE33171692143422229D319 (gx_cs_f7_bar5_is_prefetchable ), .I721D73CBB11DB0EC9DF361993F6A92EA
(gx_cs_f7_class_code ), .IE0DA0C810288CC00DF1F3AE622FFB08F (gx_cs_f7_device_id ), .IEB4CAA0AE4F26FAC1DAA6B9884179DEA
(gx_cs_f7_int_count ), .I070D33CDFCF15FB7B4DD88019C0E39E2 (gx_cs_f7_int_pin ), .I25B649490B20A1FEC9A1AA60AB0C6D5E
(gx_cs_f7_present ), .I8302D4B9F46621BBB824B1CC96E2E724 (gx_cs_f7_revision_id ), .I26BFDE09E6F548FBAC63338567411C7E
(gx_cs_f7_subsystem_id ), .I46C5269B9FB24EF04CE2CC341C288EC7 (gx_cs_subsystem_vendor_id ), .I3C9AD458B89B2FAABD743BF4E13BF421
(gx_cs_vendor_id ), .IAB32DAC10CBDBE04FD5EDBF7A576CAF9 (I51E5032D35684B1A6595F2291E95EBFD * (I96690071F3CE4794E376870D1BB87C22
/ 32)), .I394B9366718FFFBF01944193881668C1 (gx_pcie_gen2 ), .I66C185998F46A7148163982E39BCD296 (gx_tech_lib ) )
I1F30E8154B2484DAE224B45CCEF4F59C ( .ICCFB0F435B37370076102F325BC08D20 (ix_clk_125 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(ix_rst_n ), .IEE7B9D1B054F5CACBC10351FC32D7BFA (ix_pci_rsz_f0_bar0 ), .IFE8155182FD754C22D6F7FDA1F1C1174 (ix_pci_rsz_f0_bar1 ),
.ICFA3AEC9D2E8697060447D8D8EB18A80 (ix_pci_rsz_f0_bar2 ), .I81D61D198832883CFD88EB5DEB88A32B (ix_pci_rsz_f0_bar3 ),
.I1F5A786F105B576AC15A6F25EBFB89B8 (ix_pci_rsz_f0_bar4 ), .IB9B532CA44CE4054811AB748EDD0922D (ix_pci_rsz_f0_bar5 ),
.I7FE73B332A2A7E273F8EC82CC2A0A9D1 (ix_pci_rsz_f1_bar0 ), .I8C784B1A25E6B5F5402709647F921D20 (ix_pci_rsz_f1_bar1 ),
.IAFB7D4809B407BA0A70ABF120DF37844 (ix_pci_rsz_f1_bar2 ), .IA69AD6BF563BE83DB737C644B2992470 (ix_pci_rsz_f1_bar3 ),
.IBBC01C0CF0EE486327FBEB391C90772B (ix_pci_rsz_f1_bar4 ), .I147607D1A744B7E8E0F3050C499F3A23 (ix_pci_rsz_f1_bar5 ),
.IAA6C398FE19CA194DA9436764C94079A (ix_pci_rsz_f2_bar0 ), .I6375C05D4E0F58631C8731FD2B26A7F6 (ix_pci_rsz_f2_bar1 ),
.ID25293C6DC5461B1A3E61F7A7614A6D8 (ix_pci_rsz_f2_bar2 ), .I7E0B227F296E6A7FA770C68AB70324DD (ix_pci_rsz_f2_bar3 ),
.I1187CE134A1A3347BF94366BE4D44B3F (ix_pci_rsz_f2_bar4 ), .I0C7C3FDEC159F63C155144A19841E5BC (ix_pci_rsz_f2_bar5 ),
.IF0C365E1D4BC8B2941DE257EF66C8FE4 (ix_pci_rsz_f3_bar0 ), .I1646E818A90159BC4FF7AA119272C460 (ix_pci_rsz_f3_bar1 ),
.I05AD49E3884F0E62FA36DCFB88E5C22E (ix_pci_rsz_f3_bar2 ), .I348CE8EA5A014339F820FDCAFC214867 (ix_pci_rsz_f3_bar3 ),
.ICF2AC2986B60A3FD41ECFB74C4756D10 (ix_pci_rsz_f3_bar4 ), .I13B899B342E8552CACED9E20E0F5FD83 (ix_pci_rsz_f3_bar5 ),
.I068B3206EC02BBE1225E3FD649DCAC3E (ix_pci_rsz_f4_bar0 ), .I15D8A1D8934ABE732F753BC8A130129E (ix_pci_rsz_f4_bar1 ),
.IFE8F569C18FBA7444D4832F2CB5D2D69 (ix_pci_rsz_f4_bar2 ), .I51FF9F99E3F92A151FD3D6BBAAC89FB6 (ix_pci_rsz_f4_bar3 ),
.IA4118298EF0A9C92D5D3ECB07C8AE533 (ix_pci_rsz_f4_bar4 ), .I7D032A1E448C6F22898894E594BF2DD3 (ix_pci_rsz_f4_bar5 ),
.I67444F97CA6B95448FAFAE30BC1EA4A3 (ix_pci_rsz_f5_bar0 ), .ID449FF330193AAA4C7942F23F18CEF54 (ix_pci_rsz_f5_bar1 ),
.I3CABF30E4ECE3E02DF7BB2FAE8895026 (ix_pci_rsz_f5_bar2 ), .I46EAD98AAF05965858087C6CCDFEAFFD (ix_pci_rsz_f5_bar3 ),
.I1967BD95F38270D97B0A4B182C5D8F0E (ix_pci_rsz_f5_bar4 ), .ICDB8224D569BB5A5B320A26E2B451BAC (ix_pci_rsz_f5_bar5 ),
.I8220BA29B6C07A3A107C2B3234F5FB06 (ix_pci_rsz_f6_bar0 ), .I7DA2457F5006629E45D78C4FC855DCF8 (ix_pci_rsz_f6_bar1 ),
.IBB764C0D62FD349F6FB3F52A8C78424E (ix_pci_rsz_f6_bar2 ), .IE074E5B8DF895724AB3B5023BAC298BC (ix_pci_rsz_f6_bar3 ),
.IDA2FA24095F53E4EBBAC1E30772082B4 (ix_pci_rsz_f6_bar4 ), .I27FBA72EC841BBBDD25E028A08A3F06C (ix_pci_rsz_f6_bar5 ),
.I4FB68E387DB515A46DAA2DABF6E0D1D8 (ix_pci_rsz_f7_bar0 ), .IBA4DC2E68E546946B55995DB900F74F7 (ix_pci_rsz_f7_bar1 ),
.I28A9F4DDE0D0FFADF8668EFA99C6DA03 (ix_pci_rsz_f7_bar2 ), .IE02A2D602D1C83798270DD49EF6A4D23 (ix_pci_rsz_f7_bar3 ),
.I4DBB86A2215D89E37CDE4EC7DC8435C5 (ix_pci_rsz_f7_bar4 ), .I8DCB72E575B62CC266039827C0238E34 (ix_pci_rsz_f7_bar5 ),
.I8B1798242C3B0E655181D0D365813614 (I220A96CF74656D5120C8D113E4B1ED55 ), .IE145222FDBDC80109E12FA72D3D3C655 (IBE8D7D536CBDF087E7E00B93DA215E3D ),
.ID43AC1009727D128F1C5DFE4640CA5AB (I4DC446D96F0774A667A70D52D9392874 ), .IB610431939CB8180EAC2403672BAF58D (I3FF9BAFBF91288E78D7EA6DD95DB3A40 ),
.I3C7A9FA839F554D8898020C4831479E2 (IE67E5659AC07E2D371890CDACFA6ED42 ), .I74A0936EE8FD1443A2C6745A4F3F6B5E (I18137FEBF7FA4CE04FDE793386121F57 ),
.I369BA2FFB5D41DF25F9BC3AB126D6607 (I0B37325C0AB5EEA3148286371EB202D1 ), .I1C0271AD5E8E9E9164909E468AD0B212 (ix_pci_int_req ),
.I6EC1BE4B18EC6AA3D88A5D45B614565E (IFDD7175F3E1142C3A73A9731A4DF519B ), .IB907C2624CE144BCE5A772623C46F678 ({9{I026F76BAC2C8DF5D427631DEA76B062F }}),
.I3FF97406B3ED373B267711109A980AF9 (IB9BCD6E1EA621FDF5DD229996ADC5F8F ), .I24C403550AE065D7D1B7266142886226 (I026F76BAC2C8DF5D427631DEA76B062F ),
.I438B8BD876741F9B46EB770E92F808B7 (IE81C89DB2F6C737F2D82BE35AFC7DDA2 [14:0]), .I5FE75BE614D4F52DB327549B36203350
(I291FF0AF6B998FB4D8BD958CFDA1CF8C ), .I3D6C771D05CA1A769E61302C086494B8 (IEC017B3AB9F16AE871D5253A5257D941 [31:0]),
.I357B3043EDACE3EBECE8F54D79B9F90A (I87343FD56CEFDCB10F9A272CF1F0CA8E ), .I0AAD559CF33A5CBA597990658774FEB3 (IB8F3718FAD7719FD71FDE3B0DE8D7445 ),
.I923204A95D8CBB206587CF32BEDCF4EF (I678B3227DE7FFEFE726CE68123B91F8D ), .ICF9D8FD31DFC7D20DAF939C6D75F1518 (I4BA2D171F5FD7E0FEACB9DF4C87DDC19 ),
.I20CD33DEFBDF51E2A5352736B083738D (IC0197882115D001485B37646159E234E ), .IDF550B17734BF16B7E410B19BB31E276 (IB1AAAED8469CADFA3AB4BF806A8466B6 ),
.I8ED9B9C1D9F58C5D06A9443AD901E8C6 (IA6774F4F4F3AF83C6A9E233DB00F89A0 ), .IA976D63BEECA80DCE31365CF56EC0248 (IFFF50035216FD68A74F8164F0EE74689 ),
.I5E3CE5AF5C34D232BFB139B63D9912B4 (IF9A16909C25386742335A246DEDE12E8 ), .IBEF3E5F9395E2C7822AE03D6461DEBBB (I5078F81AE0F5DCD4CC2ABEE2CEF9C827 ),
.I7E6CFD6A7DCAB9CD2188D044C7D716A6 (IB55475954FE95F83F22B1C2FB76FAEC7 ), .I3A34691662384260F0524DD7F650E75A (I31980ABC07D19BA89784085C7754DE42 ),
.IC2F58AB5028C1D2C53C6EF47A4975D0A (IE1F9397E899B4E938A0D54FC51445C13 ), .I112E0A79129A8BC6DD4C13647C31F8A0 (IDE0F2D42601304C0E0CCD60778B3938F ),
.ID3E7F4B58943229FEE6313A36B3F8693 (I395C5996AD91572D0F6652373B6018E7 ), .I1FDEC1735547330C00A0B8DFE1FB10C3 (I5B507E107F91FDBF0B2EEF7DD9AE40C5 ),
.IBD6A65D48B4A68CA0D2A82F79053757B (IBAE868C7DE15BF2F751B0177B798BDCD ), .I42A419EB6EB8D11234AC3B2BCA0AE593 (IAF2A92B584FD036A9F751EB8F3FA7ACD ),
.IA41AC3CC6BC050DDC172724AB311315B (I5CF35907FA895D81AAC1AAFED86DBE1F ), .I31CF69FF368B36B4D6612DF16B3ABC6B (I1BAAE01807D45E9F21D2ACB2BCB4F621 ),
.I439AF6D496491F5F7C23217209B43C31 (ID872B1CCC580E5915A782E136C7A691B ), .IFE4A8CBA73734C6F0F0A078027E053D4 (IFFB9EED620356BDFB94697DB3606174F ),
.ID7A2A8B1E9D92B60194D5FAFAAB15208 (I2C072E656BFCADF4877B42244D6D2307 ), .IF274FAF97F5BACD693913BB418717A9D (IB96A9322FAF5941DF70737CA69F152A3 ),
.I270ED686C2EF2C1C8B5B55EC4A5AAE84 (I9625E96E33563830A2A0ED7263124B10 ), .ID5CCD4858CB5CC1B2EDEC682C7DE5AAD (I1B43D1CE930FCA067FA31726F2C15FEE ),
.I7D901091F9E0741061C75B54467D48A0 (I697639B04C0F4B6F9764F8122329FB7C ) ); I7639B3DE6448BF04A6DF404C0FEDBA75 # (
.I7292F55C07BFD7FB8A60D29FFC186275 (I96690071F3CE4794E376870D1BB87C22 ), .IDB751C3DD512B8355CF27001F983880A (gx_ipx_data_sz ),
.I99651B9F47529E0ADC5349B57C84E531 (I90D984439DDA58639C67AC709C0E6CC9 ), .ICED1C5B792370B25488CFA18FE5E472E (I31F00D08C3CE05C5A25E18130CAFEAD5 ),
.I0AEF008AE3BC7E23C49F86BC2B344750 (I51E5032D35684B1A6595F2291E95EBFD ), .I026FA76AB836F95856A0F400EDF284FA (IF3D376C350B88011F1FC2F939263D178 ),
.I66C185998F46A7148163982E39BCD296 (gx_tech_lib ), .I6684631E4DAAC3FB7551EF267A7E3D73 (gx_wbm_data_sz ), .I3A59A966031A54015DBF77A68A5A82D3
(gx_wbs_data_sz ) ) I50AE61DF7EF91EA9267CD28222E12D54 ( .ICCFB0F435B37370076102F325BC08D20 (ix_clk_125 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(ix_rst_n ), .I488999E90FEFB5E25518723EB6105532 (ix_ipx_tx_ca_cpld ), .IB064E00468F70C38840D1D271524C6C8 (ix_ipx_tx_ca_cplh ),
.IE4E19EA6F3F828B3B44ED1E4D36558F7 (ix_ipx_tx_ca_npd ), .I537C738B170D60A42A1F6FDA4547BACC (ix_ipx_tx_ca_nph ),
.IA29842BA67669CD8D75483E633C363F0 (ix_ipx_tx_ca_pd ), .IB9E3BDBEE7C442BA69CD12711DA40F71 (ix_ipx_tx_ca_ph ), .IABD5FBD9A9966396ACABECC997D287C6
(ix_ipx_tx_rdy ), .IFCFFF8448F5E6821B40C6CEE3548693A (ix_ipx_tx_val ), .I5CE5D2469FD5560C1773C754FC1E0C4A (ix_ipx_pcie_linkw ),
.ID965E2D89D1047516134A3EED50CB8AE (ix_ipx_pcie_rate ), .I884F4ADE09FABBA20600F67BC1A50FE7 (I6609F40DB9BF2AAD262974646AD5EBE5 ),
.I61E8E6981294A3342BDF5596043A2DFA (IAE96F702FDFFAF4D7DD2303A7E5CAA82 ), .I2F5C52C0CABA5EFAF34A96BC39DA8F96 (I314F20E260B367A911975FFD9E094426 ),
.I0BA940AC86B853EFCE63667C128E2DF4 (IE5A769A04E820A9426CF9BB3B0A13E3C ), .ID176017A6F96653AFD707B70D22BEA8C (IF35E88F0598148E05EAD3AB0F7ED2F9E ),
.IE8C34BE7792A66A23CB1C7A5CFF55BBF (I7A68BADCCB87652618C1488B18D4A938 ), .IA5896E672427191F9A0B4ED1C9301313 (IFFB9EED620356BDFB94697DB3606174F ),
.I0317313DEECD8AC19E98BA2F1C27E0A9 (I2C072E656BFCADF4877B42244D6D2307 ), .IFDB2ACAC637F40CDDFBB20A3AFD9A401 (IB96A9322FAF5941DF70737CA69F152A3 ),
.IE4C3654339F6BF285840C2AB868371A1 (I10A77B5F026A0F0CC0D1B6C8CD9C0746 ), .I5F40D6DD3270B21E2E90925F127E6477 (I5257580F4980618A2A58EA7899EEC7B5 ),
.I33A8C146E90D24E54E605500849CD461 (ICBA9D9788BB5A0277607D0E038FE4333 ), .I42D2723FE4CDE4AF565DD01BD32BB8AC (I4A399AD6EACAD372F1F0ED553AF29E10 ),
.I8E99DEF5C63C6A55606BD30E4BE8E3FB (ICCEE7A1D3C2702A0766B02D0E4CD1F5A ), .IC3760F6E74F9AA61561390CC1466FC1A (I9625E96E33563830A2A0ED7263124B10 ),
.I582940C94DBA710A62923187D833E8E6 (ID0B88392A9310E618D259D3AE74555DF ), .IDFCF1C6E3889548A5224E9568D7E2E22 (I11AAD529B8C632E2B3F7E5810F154FAE ),
.I241490D6913C41E3972F651398E36880 (I6E8F4533B895189C22AD2D5F06D2C022 ), .IA127FE276B1C05C6A690F8454BBF510B (IB9BCD6E1EA621FDF5DD229996ADC5F8F ),
.I0ED116F3061ADCE682AE68F0A5003CBF (I6037B76B56AF44132A3D98CA48DE55B0 ), .IB33B8D629A269D1BC3D79902EE2EB312 (I9A5D7FA3649743F4C12D7A2A0F5D00B9 ),
.I1E494BBA2ECB063404DBB73667CC7E8D (IB72EDE3F33BC320C4BB54A891CA0124E ), .I4A4976CAF016EA789DCDB7AA131246C3 (I597BFE708F080A1AC7F68B18B2D32AEF ),
.I5ADFC7E7F8B570F5258C2813D0020950 (I452B7C3155C15AA425E22E8ACF0B4BDF ), .I1FD27F5D298FA5493F3F510610F19E4E (IBCEC5B979CD682F2C507E946AAC6F86F ),
.IAFF3235BDF22DE6B7D7DBF12451FA2FE (I443AE8A2A80F3D4BC5B0F9739DC268B7 ), .I5FFD1878342C11E50C1617928EBB38D7 (IF35D2DA8FDBB83C8C227111A766BE7D7 ),
.I27766E6DFBDE7E37CDB16F4E2C0E1DD4 (I026F76BAC2C8DF5D427631DEA76B062F ), .I520751EAD225B5BFC3D7E0ACB7BC6405 (IE9523C108AFE8D1C07903BFCE449B9F8 )
); credit_config IE31D1703EF68AF964E0E8781D43B7506 ( .ox_fc_cpld_infinite ( ), .ox_fc_cplh_infinite ( ), .ox_fc_npd_infinite
(IFD9B46ACBF1F17D2A8C784B3B4B2901E ), .ox_fc_nph_infinite (I42C3C6068A9CD9CB33558F95CD336652 ), .ox_fc_pd_infinite
(I39F7612EB75C5A11AF508BF344CD51B8 ), .ox_fc_ph_infinite (ICF4A96ABEB44A00DC9123A0C152DC218 ), .ox_io_space_sel
( ), .ox_hw_rev ( ), .ox_subsys_id ( ) ); I35D01845B6D15D59E4E7B95EDE6F3368 #( .I7292F55C07BFD7FB8A60D29FFC186275
(IEF532EA44160288B0ED6812C670E4CDB ), .IB71844FFA3AB85FEF45EAB4D35395752 (IF3D376C350B88011F1FC2F939263D178 ), .IDB9D60794264C5F8E5363941194A797B
(gx_nr_wb_tgts ), .I66C185998F46A7148163982E39BCD296 (gx_tech_lib ), .ID7C7F9F2E39BEBEE2ACFA8040034E48D (gx_wbm_adr_sz )
) IF18997A3ADD4120C792F1288A675E468 ( .ICCFB0F435B37370076102F325BC08D20 (ix_clk_125 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(ix_rst_n ), .IF87783FDF111A8E49EAC36F1DDFCBA80 (ix_wbm_ack ), .IF9D5978BE23690B1D4D13EF2AD676C6F (ix_wbm_dat ),
.IDC6EA54AB52AEAD439CEF7521615AE1B (IE81C89DB2F6C737F2D82BE35AFC7DDA2 ), .I6ED49B5BED4BA586759FFDCC7B3B7FF8 (I599F86FA1B9AEED5B32EE8B27DFFFACE ),
.I8E2F7CF6E50B95A483351A1836EB23AC (IDCB78AD56EF8FEF35AAF4DED8D1F87B6 ), .I506D2FCB600E0189274870B654E65B64 (IEC017B3AB9F16AE871D5253A5257D941 ),
.I141300E29D7EF4A0D8B71CB7469A7B90 (IB8F3718FAD7719FD71FDE3B0DE8D7445 ), .I9AF8DD3F367CE82DF45437DB546EAAD3 (I5EB48F61C7554EB021FC36EC1077B4B1 ),
.I42D281FF99DC79A9AD9E7DF0AEB073A7 (I7681E0E609A03559F13166ACF7852905 ), .I3068B33EE97A971AE7F0CF17705AA6DC (I507A0A1A3C69E79845F5C15AFFAF6595 ),
.IFCBA19703D55B4610B3F4174C5B8833A (IDB0B420EA96A60B402FECD3AE3620DCC ), .IC3CC91D317012C130AC9E2A126F71C64 (I678B3227DE7FFEFE726CE68123B91F8D ),
.I561BE0F01153FC1AADDEB08B34B545B6 (I6C86D46877E4F106568E7404A48B3614 ), .IB86AF6EBEEA3CE1BF22AE1AF7CC8481F (I1EBAB68345C1F3BB0BA0E7EF6A0A1648 ),
.I94E3D00BBC13BF182097A25D63288C2C (I25EB4135E1552B388D1686480F82F884 ), .I8B25F4450817FC10E1E3DC6B500C9F5A (IECA17FE57E485E6400F2DB42821DD251 ),
.I26C902CE18647F75561AD003E260B048 (I02736097A9414A8EE96C59AC2C4D85D6 ), .IA5CEBFC654EDCA4107594F388D5BC88A (IE7216A06BFCE79862D756B0F69D722FB ),
.I27627079DD78A85D26D85DC0C53D835F (I109964893AEF92F63170615855D13B10 ), .I0205131FB84BB0F9F8AD5CC00E5E861D (I2407989C7097E49E194FF778C1BA69FD ),
.IDA581E8478C8224118EF4E6B8EE8DDFE (IFDE36B1D5ECEDDC8E1D64BAC3AB778F5 ), .IA36C0DD0DE88B03FA61EF35103D22DF0 (IF61A4C9125864F891B9412F7F8A38722 )
); ID81B7D29F9F1B2882EE754B639B67517 #( .I7292F55C07BFD7FB8A60D29FFC186275 (gx_wbs_data_sz ), .IC3CEA40E2663BA267FBD739EE37AFBE9
(I31F00D08C3CE05C5A25E18130CAFEAD5 * (I96690071F3CE4794E376870D1BB87C22 / gx_wbm_data_sz )), .IAB32DAC10CBDBE04FD5EDBF7A576CAF9
(IF3D376C350B88011F1FC2F939263D178 * (I96690071F3CE4794E376870D1BB87C22 / gx_wbm_data_sz )), .IB941270487D75F8FAA82F3DF028B6FC6
(I96690071F3CE4794E376870D1BB87C22 ), .IFB129920FFBFCFD17ADB3180F882E8E1 (gx_wbs_adr_sz ), .I66C185998F46A7148163982E39BCD296
(gx_tech_lib ) ) I55AD3DB98631F7D24697571C1AE7D521 ( .ICCFB0F435B37370076102F325BC08D20 (ix_clk_125 ), .I9ED2A9117D3AEAF54CBA7AD69083BCB7
(ix_rst_n ), .IC680604FB338D55088F12313CDF2B03E (I4BA2D171F5FD7E0FEACB9DF4C87DDC19 ), .IF17B1273FDE2637DBFCD3D142F80E5D5
(I395C5996AD91572D0F6652373B6018E7 ), .I44E00CA48D123AE945CB7C612A95BFE6 (I5B507E107F91FDBF0B2EEF7DD9AE40C5 ), .I6D124B4E6D5F74B43E94949DE1CF46AA
(IAF2A92B584FD036A9F751EB8F3FA7ACD ), .I5C266315A3CF63C3FE988BB363C59AA1 (I5CF35907FA895D81AAC1AAFED86DBE1F ), .I3EEFAC16E2400143CD0547F03531871C
(IB552918C70C5F8374FC906E0C2225F89 ), .I77DB6FE5680F7C0F4CCBA7F787115DDC (IE593D61A89622FBF1D4D61DBF77B0759 ), .I7AC0939DFAAFF38545186E63551C4452
(I25B75CE7CA22EBCC6B686F9FD442035C ), .I10E4ABD5838C4A0B5C07B5A66417237D (I6E8F4533B895189C22AD2D5F06D2C022 ), .I3FF97406B3ED373B267711109A980AF9
(I6037B76B56AF44132A3D98CA48DE55B0 ), .I238A13C6F03704581F9A0A170F852FB4 (IF35D2DA8FDBB83C8C227111A766BE7D7 ), .I24C403550AE065D7D1B7266142886226
(IE9523C108AFE8D1C07903BFCE449B9F8 ), .IDC6EA54AB52AEAD439CEF7521615AE1B (ix_wbs_adr ), .IC93EB5988EC451F72626A919FE396C61
(ix_wbs_bte ), .I6ED49B5BED4BA586759FFDCC7B3B7FF8 (ix_wbs_cti ), .I8E2F7CF6E50B95A483351A1836EB23AC (ix_wbs_cyc ),
.I506D2FCB600E0189274870B654E65B64 (ix_wbs_dat ), .I1304D1B0EBC59FFD53EF6CD7A8537E4D (ix_wbs_sel ), .I141300E29D7EF4A0D8B71CB7469A7B90
(ix_wbs_stb ), .IC3CC91D317012C130AC9E2A126F71C64 (ix_wbs_we ), .I7244B3A041E4EF91034ED304D36B4585 (IFDD7175F3E1142C3A73A9731A4DF519B ),
.IC3E8DB22A270F4E2527F04E7E81EFA46 (IF35E88F0598148E05EAD3AB0F7ED2F9E ), .IAEC671D12B80E2CC6E3D591A98E27230 (I7A68BADCCB87652618C1488B18D4A938 ),
.IA449B4CEADDC750F5446E3B900C14AA4 (IE5A769A04E820A9426CF9BB3B0A13E3C ), .IFA413F55A4E38AA4A08DC60DCCB7553D (I5257580F4980618A2A58EA7899EEC7B5 ),
.I80F26623B387879BCA3F00C252D0129E (ICBA9D9788BB5A0277607D0E038FE4333 ), .IFC7E490A5AF630CDD63895FB063ABE29 (I10A77B5F026A0F0CC0D1B6C8CD9C0746 ),
.IEBE9989B3828CC1007CD10E6FBB2E76C (ICCEE7A1D3C2702A0766B02D0E4CD1F5A ), .I270ED686C2EF2C1C8B5B55EC4A5AAE84 (ID0B88392A9310E618D259D3AE74555DF ),
.IDA581E8478C8224118EF4E6B8EE8DDFE (IAB567E212EF35BD2AA033B83F2307D63 ), .I197028CF3B48BF15266050E66E13618E (IC3E05B0E9AC8F202F65F1764031827B8 )
); endmodule 
